magic
tech sky130A
magscale 1 2
timestamp 1679496889
<< obsli1 >>
rect 1104 2159 102856 101745
<< obsm1 >>
rect 14 2128 103210 102264
<< metal2 >>
rect 18 103200 74 104000
rect 662 103200 718 104000
rect 1306 103200 1362 104000
rect 1950 103200 2006 104000
rect 2594 103200 2650 104000
rect 3238 103200 3294 104000
rect 3882 103200 3938 104000
rect 4526 103200 4582 104000
rect 5170 103200 5226 104000
rect 5814 103200 5870 104000
rect 6458 103200 6514 104000
rect 7746 103200 7802 104000
rect 8390 103200 8446 104000
rect 9034 103200 9090 104000
rect 9678 103200 9734 104000
rect 10322 103200 10378 104000
rect 10966 103200 11022 104000
rect 11610 103200 11666 104000
rect 12254 103200 12310 104000
rect 12898 103200 12954 104000
rect 13542 103200 13598 104000
rect 14186 103200 14242 104000
rect 14830 103200 14886 104000
rect 15474 103200 15530 104000
rect 16118 103200 16174 104000
rect 16762 103200 16818 104000
rect 17406 103200 17462 104000
rect 18050 103200 18106 104000
rect 18694 103200 18750 104000
rect 19338 103200 19394 104000
rect 19982 103200 20038 104000
rect 20626 103200 20682 104000
rect 21270 103200 21326 104000
rect 21914 103200 21970 104000
rect 22558 103200 22614 104000
rect 23202 103200 23258 104000
rect 23846 103200 23902 104000
rect 25134 103200 25190 104000
rect 25778 103200 25834 104000
rect 26422 103200 26478 104000
rect 27066 103200 27122 104000
rect 27710 103200 27766 104000
rect 28354 103200 28410 104000
rect 28998 103200 29054 104000
rect 29642 103200 29698 104000
rect 30286 103200 30342 104000
rect 30930 103200 30986 104000
rect 31574 103200 31630 104000
rect 32218 103200 32274 104000
rect 32862 103200 32918 104000
rect 33506 103200 33562 104000
rect 34150 103200 34206 104000
rect 34794 103200 34850 104000
rect 35438 103200 35494 104000
rect 36082 103200 36138 104000
rect 36726 103200 36782 104000
rect 37370 103200 37426 104000
rect 38014 103200 38070 104000
rect 38658 103200 38714 104000
rect 39302 103200 39358 104000
rect 39946 103200 40002 104000
rect 40590 103200 40646 104000
rect 41234 103200 41290 104000
rect 41878 103200 41934 104000
rect 43166 103200 43222 104000
rect 43810 103200 43866 104000
rect 44454 103200 44510 104000
rect 45098 103200 45154 104000
rect 45742 103200 45798 104000
rect 46386 103200 46442 104000
rect 47030 103200 47086 104000
rect 47674 103200 47730 104000
rect 48318 103200 48374 104000
rect 48962 103200 49018 104000
rect 49606 103200 49662 104000
rect 50250 103200 50306 104000
rect 50894 103200 50950 104000
rect 51538 103200 51594 104000
rect 52182 103200 52238 104000
rect 52826 103200 52882 104000
rect 53470 103200 53526 104000
rect 54114 103200 54170 104000
rect 54758 103200 54814 104000
rect 55402 103200 55458 104000
rect 56046 103200 56102 104000
rect 56690 103200 56746 104000
rect 57334 103200 57390 104000
rect 57978 103200 58034 104000
rect 58622 103200 58678 104000
rect 59266 103200 59322 104000
rect 60554 103200 60610 104000
rect 61198 103200 61254 104000
rect 61842 103200 61898 104000
rect 62486 103200 62542 104000
rect 63130 103200 63186 104000
rect 63774 103200 63830 104000
rect 64418 103200 64474 104000
rect 65062 103200 65118 104000
rect 65706 103200 65762 104000
rect 66350 103200 66406 104000
rect 66994 103200 67050 104000
rect 67638 103200 67694 104000
rect 68282 103200 68338 104000
rect 68926 103200 68982 104000
rect 69570 103200 69626 104000
rect 70214 103200 70270 104000
rect 70858 103200 70914 104000
rect 71502 103200 71558 104000
rect 72146 103200 72202 104000
rect 72790 103200 72846 104000
rect 73434 103200 73490 104000
rect 74078 103200 74134 104000
rect 74722 103200 74778 104000
rect 75366 103200 75422 104000
rect 76010 103200 76066 104000
rect 76654 103200 76710 104000
rect 77942 103200 77998 104000
rect 78586 103200 78642 104000
rect 79230 103200 79286 104000
rect 79874 103200 79930 104000
rect 80518 103200 80574 104000
rect 81162 103200 81218 104000
rect 81806 103200 81862 104000
rect 82450 103200 82506 104000
rect 83094 103200 83150 104000
rect 83738 103200 83794 104000
rect 84382 103200 84438 104000
rect 85026 103200 85082 104000
rect 85670 103200 85726 104000
rect 86314 103200 86370 104000
rect 86958 103200 87014 104000
rect 87602 103200 87658 104000
rect 88246 103200 88302 104000
rect 88890 103200 88946 104000
rect 89534 103200 89590 104000
rect 90178 103200 90234 104000
rect 90822 103200 90878 104000
rect 91466 103200 91522 104000
rect 92110 103200 92166 104000
rect 92754 103200 92810 104000
rect 93398 103200 93454 104000
rect 94042 103200 94098 104000
rect 94686 103200 94742 104000
rect 95974 103200 96030 104000
rect 96618 103200 96674 104000
rect 97262 103200 97318 104000
rect 97906 103200 97962 104000
rect 98550 103200 98606 104000
rect 99194 103200 99250 104000
rect 99838 103200 99894 104000
rect 100482 103200 100538 104000
rect 101126 103200 101182 104000
rect 101770 103200 101826 104000
rect 102414 103200 102470 104000
rect 103058 103200 103114 104000
rect 103702 103200 103758 104000
rect 4208 2128 4528 101776
rect 4868 2128 5188 101776
rect 5528 2128 5848 101776
rect 6188 2128 6508 101776
rect 34928 2128 35248 101776
rect 35588 2128 35908 101776
rect 36248 2128 36568 101776
rect 36908 2128 37228 101776
rect 65648 2128 65968 101776
rect 66308 2128 66628 101776
rect 66968 2128 67288 101776
rect 67628 2128 67948 101776
rect 96368 2128 96688 101776
rect 97028 2128 97348 101776
rect 97688 2128 98008 101776
rect 98348 2128 98668 101776
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103702 0 103758 800
<< obsm2 >>
rect 130 103144 606 103465
rect 774 103144 1250 103465
rect 1418 103144 1894 103465
rect 2062 103144 2538 103465
rect 2706 103144 3182 103465
rect 3350 103144 3826 103465
rect 3994 103144 4470 103465
rect 4638 103144 5114 103465
rect 5282 103144 5758 103465
rect 5926 103144 6402 103465
rect 6570 103144 7690 103465
rect 7858 103144 8334 103465
rect 8502 103144 8978 103465
rect 9146 103144 9622 103465
rect 9790 103144 10266 103465
rect 10434 103144 10910 103465
rect 11078 103144 11554 103465
rect 11722 103144 12198 103465
rect 12366 103144 12842 103465
rect 13010 103144 13486 103465
rect 13654 103144 14130 103465
rect 14298 103144 14774 103465
rect 14942 103144 15418 103465
rect 15586 103144 16062 103465
rect 16230 103144 16706 103465
rect 16874 103144 17350 103465
rect 17518 103144 17994 103465
rect 18162 103144 18638 103465
rect 18806 103144 19282 103465
rect 19450 103144 19926 103465
rect 20094 103144 20570 103465
rect 20738 103144 21214 103465
rect 21382 103144 21858 103465
rect 22026 103144 22502 103465
rect 22670 103144 23146 103465
rect 23314 103144 23790 103465
rect 23958 103144 25078 103465
rect 25246 103144 25722 103465
rect 25890 103144 26366 103465
rect 26534 103144 27010 103465
rect 27178 103144 27654 103465
rect 27822 103144 28298 103465
rect 28466 103144 28942 103465
rect 29110 103144 29586 103465
rect 29754 103144 30230 103465
rect 30398 103144 30874 103465
rect 31042 103144 31518 103465
rect 31686 103144 32162 103465
rect 32330 103144 32806 103465
rect 32974 103144 33450 103465
rect 33618 103144 34094 103465
rect 34262 103144 34738 103465
rect 34906 103144 35382 103465
rect 35550 103144 36026 103465
rect 36194 103144 36670 103465
rect 36838 103144 37314 103465
rect 37482 103144 37958 103465
rect 38126 103144 38602 103465
rect 38770 103144 39246 103465
rect 39414 103144 39890 103465
rect 40058 103144 40534 103465
rect 40702 103144 41178 103465
rect 41346 103144 41822 103465
rect 41990 103144 43110 103465
rect 43278 103144 43754 103465
rect 43922 103144 44398 103465
rect 44566 103144 45042 103465
rect 45210 103144 45686 103465
rect 45854 103144 46330 103465
rect 46498 103144 46974 103465
rect 47142 103144 47618 103465
rect 47786 103144 48262 103465
rect 48430 103144 48906 103465
rect 49074 103144 49550 103465
rect 49718 103144 50194 103465
rect 50362 103144 50838 103465
rect 51006 103144 51482 103465
rect 51650 103144 52126 103465
rect 52294 103144 52770 103465
rect 52938 103144 53414 103465
rect 53582 103144 54058 103465
rect 54226 103144 54702 103465
rect 54870 103144 55346 103465
rect 55514 103144 55990 103465
rect 56158 103144 56634 103465
rect 56802 103144 57278 103465
rect 57446 103144 57922 103465
rect 58090 103144 58566 103465
rect 58734 103144 59210 103465
rect 59378 103144 60498 103465
rect 60666 103144 61142 103465
rect 61310 103144 61786 103465
rect 61954 103144 62430 103465
rect 62598 103144 63074 103465
rect 63242 103144 63718 103465
rect 63886 103144 64362 103465
rect 64530 103144 65006 103465
rect 65174 103144 65650 103465
rect 65818 103144 66294 103465
rect 66462 103144 66938 103465
rect 67106 103144 67582 103465
rect 67750 103144 68226 103465
rect 68394 103144 68870 103465
rect 69038 103144 69514 103465
rect 69682 103144 70158 103465
rect 70326 103144 70802 103465
rect 70970 103144 71446 103465
rect 71614 103144 72090 103465
rect 72258 103144 72734 103465
rect 72902 103144 73378 103465
rect 73546 103144 74022 103465
rect 74190 103144 74666 103465
rect 74834 103144 75310 103465
rect 75478 103144 75954 103465
rect 76122 103144 76598 103465
rect 76766 103144 77886 103465
rect 78054 103144 78530 103465
rect 78698 103144 79174 103465
rect 79342 103144 79818 103465
rect 79986 103144 80462 103465
rect 80630 103144 81106 103465
rect 81274 103144 81750 103465
rect 81918 103144 82394 103465
rect 82562 103144 83038 103465
rect 83206 103144 83682 103465
rect 83850 103144 84326 103465
rect 84494 103144 84970 103465
rect 85138 103144 85614 103465
rect 85782 103144 86258 103465
rect 86426 103144 86902 103465
rect 87070 103144 87546 103465
rect 87714 103144 88190 103465
rect 88358 103144 88834 103465
rect 89002 103144 89478 103465
rect 89646 103144 90122 103465
rect 90290 103144 90766 103465
rect 90934 103144 91410 103465
rect 91578 103144 92054 103465
rect 92222 103144 92698 103465
rect 92866 103144 93342 103465
rect 93510 103144 93986 103465
rect 94154 103144 94630 103465
rect 94798 103144 95918 103465
rect 96086 103144 96562 103465
rect 96730 103144 97206 103465
rect 97374 103144 97850 103465
rect 98018 103144 98494 103465
rect 98662 103144 99138 103465
rect 99306 103144 99782 103465
rect 99950 103144 100426 103465
rect 100594 103144 101070 103465
rect 101238 103144 101714 103465
rect 101882 103144 102358 103465
rect 102526 103144 103002 103465
rect 103170 103144 103204 103465
rect 20 101832 103204 103144
rect 20 2072 4152 101832
rect 4584 2072 4812 101832
rect 5244 2072 5472 101832
rect 5904 2072 6132 101832
rect 6564 2072 34872 101832
rect 35304 2072 35532 101832
rect 35964 2072 36192 101832
rect 36624 2072 36852 101832
rect 37284 2072 65592 101832
rect 66024 2072 66252 101832
rect 66684 2072 66912 101832
rect 67344 2072 67572 101832
rect 68004 2072 96312 101832
rect 96744 2072 96972 101832
rect 97404 2072 97632 101832
rect 98064 2072 98292 101832
rect 98724 2072 103204 101832
rect 20 856 103204 2072
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 14774 856
rect 14942 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21214 856
rect 21382 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30230 856
rect 30398 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34094 856
rect 34262 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37314 856
rect 37482 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39246 856
rect 39414 31 39890 856
rect 40058 31 40534 856
rect 40702 31 41178 856
rect 41346 31 41822 856
rect 41990 31 42466 856
rect 42634 31 43110 856
rect 43278 31 43754 856
rect 43922 31 44398 856
rect 44566 31 45042 856
rect 45210 31 45686 856
rect 45854 31 46330 856
rect 46498 31 46974 856
rect 47142 31 47618 856
rect 47786 31 48262 856
rect 48430 31 48906 856
rect 49074 31 49550 856
rect 49718 31 50194 856
rect 50362 31 50838 856
rect 51006 31 51482 856
rect 51650 31 52126 856
rect 52294 31 53414 856
rect 53582 31 54058 856
rect 54226 31 54702 856
rect 54870 31 55346 856
rect 55514 31 55990 856
rect 56158 31 56634 856
rect 56802 31 57278 856
rect 57446 31 57922 856
rect 58090 31 58566 856
rect 58734 31 59210 856
rect 59378 31 59854 856
rect 60022 31 60498 856
rect 60666 31 61142 856
rect 61310 31 61786 856
rect 61954 31 62430 856
rect 62598 31 63074 856
rect 63242 31 63718 856
rect 63886 31 64362 856
rect 64530 31 65006 856
rect 65174 31 65650 856
rect 65818 31 66294 856
rect 66462 31 66938 856
rect 67106 31 67582 856
rect 67750 31 68226 856
rect 68394 31 68870 856
rect 69038 31 69514 856
rect 69682 31 70802 856
rect 70970 31 71446 856
rect 71614 31 72090 856
rect 72258 31 72734 856
rect 72902 31 73378 856
rect 73546 31 74022 856
rect 74190 31 74666 856
rect 74834 31 75310 856
rect 75478 31 75954 856
rect 76122 31 76598 856
rect 76766 31 77242 856
rect 77410 31 77886 856
rect 78054 31 78530 856
rect 78698 31 79174 856
rect 79342 31 79818 856
rect 79986 31 80462 856
rect 80630 31 81106 856
rect 81274 31 81750 856
rect 81918 31 82394 856
rect 82562 31 83038 856
rect 83206 31 83682 856
rect 83850 31 84326 856
rect 84494 31 84970 856
rect 85138 31 85614 856
rect 85782 31 86258 856
rect 86426 31 86902 856
rect 87070 31 88190 856
rect 88358 31 88834 856
rect 89002 31 89478 856
rect 89646 31 90122 856
rect 90290 31 90766 856
rect 90934 31 91410 856
rect 91578 31 92054 856
rect 92222 31 92698 856
rect 92866 31 93342 856
rect 93510 31 93986 856
rect 94154 31 94630 856
rect 94798 31 95274 856
rect 95442 31 95918 856
rect 96086 31 96562 856
rect 96730 31 97206 856
rect 97374 31 97850 856
rect 98018 31 98494 856
rect 98662 31 99138 856
rect 99306 31 99782 856
rect 99950 31 100426 856
rect 100594 31 101070 856
rect 101238 31 101714 856
rect 101882 31 102358 856
rect 102526 31 103002 856
rect 103170 31 103204 856
<< metal3 >>
rect 0 103368 800 103488
rect 103200 103368 104000 103488
rect 0 102688 800 102808
rect 103200 102688 104000 102808
rect 0 102008 800 102128
rect 103200 102008 104000 102128
rect 0 101328 800 101448
rect 103200 101328 104000 101448
rect 0 100648 800 100768
rect 103200 100648 104000 100768
rect 0 99968 800 100088
rect 103200 99968 104000 100088
rect 0 99288 800 99408
rect 103200 99288 104000 99408
rect 0 98608 800 98728
rect 103200 98608 104000 98728
rect 0 97928 800 98048
rect 103200 97928 104000 98048
rect 0 97248 800 97368
rect 103200 97248 104000 97368
rect 0 96568 800 96688
rect 103200 96568 104000 96688
rect 0 95888 800 96008
rect 103200 95888 104000 96008
rect 0 95208 800 95328
rect 103200 95208 104000 95328
rect 0 94528 800 94648
rect 0 93848 800 93968
rect 103200 93848 104000 93968
rect 0 93168 800 93288
rect 103200 93168 104000 93288
rect 103200 92488 104000 92608
rect 0 91808 800 91928
rect 103200 91808 104000 91928
rect 0 91128 800 91248
rect 103200 91128 104000 91248
rect 0 90448 800 90568
rect 103200 90448 104000 90568
rect 0 89768 800 89888
rect 103200 89768 104000 89888
rect 0 89088 800 89208
rect 103200 89088 104000 89208
rect 0 88408 800 88528
rect 103200 88408 104000 88528
rect 0 87728 800 87848
rect 103200 87728 104000 87848
rect 0 87048 800 87168
rect 103200 87048 104000 87168
rect 0 86368 800 86488
rect 103200 86368 104000 86488
rect 0 85688 800 85808
rect 103200 85688 104000 85808
rect 0 85008 800 85128
rect 103200 85008 104000 85128
rect 0 84328 800 84448
rect 103200 84328 104000 84448
rect 0 83648 800 83768
rect 103200 83648 104000 83768
rect 0 82968 800 83088
rect 103200 82968 104000 83088
rect 0 82288 800 82408
rect 103200 82288 104000 82408
rect 0 81608 800 81728
rect 103200 81608 104000 81728
rect 0 80928 800 81048
rect 103200 80928 104000 81048
rect 0 80248 800 80368
rect 103200 80248 104000 80368
rect 0 79568 800 79688
rect 103200 79568 104000 79688
rect 0 78888 800 79008
rect 103200 78888 104000 79008
rect 0 78208 800 78328
rect 103200 78208 104000 78328
rect 0 77528 800 77648
rect 103200 77528 104000 77648
rect 0 76848 800 76968
rect 103200 76848 104000 76968
rect 0 76168 800 76288
rect 103200 76168 104000 76288
rect 0 75488 800 75608
rect 0 74808 800 74928
rect 103200 74808 104000 74928
rect 103200 74128 104000 74248
rect 0 73448 800 73568
rect 103200 73448 104000 73568
rect 0 72768 800 72888
rect 103200 72768 104000 72888
rect 0 72088 800 72208
rect 103200 72088 104000 72208
rect 0 71408 800 71528
rect 103200 71408 104000 71528
rect 0 70728 800 70848
rect 103200 70728 104000 70848
rect 0 70048 800 70168
rect 103200 70048 104000 70168
rect 0 69368 800 69488
rect 103200 69368 104000 69488
rect 0 68688 800 68808
rect 103200 68688 104000 68808
rect 0 68008 800 68128
rect 103200 68008 104000 68128
rect 0 67328 800 67448
rect 103200 67328 104000 67448
rect 0 66648 800 66768
rect 103200 66648 104000 66768
rect 0 65968 800 66088
rect 103200 65968 104000 66088
rect 0 65288 800 65408
rect 103200 65288 104000 65408
rect 0 64608 800 64728
rect 103200 64608 104000 64728
rect 0 63928 800 64048
rect 103200 63928 104000 64048
rect 0 63248 800 63368
rect 103200 63248 104000 63368
rect 0 62568 800 62688
rect 103200 62568 104000 62688
rect 0 61888 800 62008
rect 103200 61888 104000 62008
rect 0 61208 800 61328
rect 103200 61208 104000 61328
rect 0 60528 800 60648
rect 103200 60528 104000 60648
rect 0 59848 800 59968
rect 103200 59848 104000 59968
rect 0 59168 800 59288
rect 103200 59168 104000 59288
rect 0 58488 800 58608
rect 103200 58488 104000 58608
rect 0 57808 800 57928
rect 103200 57808 104000 57928
rect 0 57128 800 57248
rect 0 56448 800 56568
rect 103200 56448 104000 56568
rect 103200 55768 104000 55888
rect 0 55088 800 55208
rect 103200 55088 104000 55208
rect 0 54408 800 54528
rect 103200 54408 104000 54528
rect 0 53728 800 53848
rect 103200 53728 104000 53848
rect 0 53048 800 53168
rect 103200 53048 104000 53168
rect 0 52368 800 52488
rect 103200 52368 104000 52488
rect 0 51688 800 51808
rect 103200 51688 104000 51808
rect 0 51008 800 51128
rect 103200 51008 104000 51128
rect 0 50328 800 50448
rect 103200 50328 104000 50448
rect 0 49648 800 49768
rect 103200 49648 104000 49768
rect 0 48968 800 49088
rect 103200 48968 104000 49088
rect 0 48288 800 48408
rect 103200 48288 104000 48408
rect 0 47608 800 47728
rect 103200 47608 104000 47728
rect 0 46928 800 47048
rect 103200 46928 104000 47048
rect 0 46248 800 46368
rect 103200 46248 104000 46368
rect 0 45568 800 45688
rect 103200 45568 104000 45688
rect 0 44888 800 45008
rect 103200 44888 104000 45008
rect 0 44208 800 44328
rect 103200 44208 104000 44328
rect 0 43528 800 43648
rect 103200 43528 104000 43648
rect 0 42848 800 42968
rect 103200 42848 104000 42968
rect 0 42168 800 42288
rect 103200 42168 104000 42288
rect 0 41488 800 41608
rect 103200 41488 104000 41608
rect 0 40808 800 40928
rect 103200 40808 104000 40928
rect 0 40128 800 40248
rect 103200 40128 104000 40248
rect 0 39448 800 39568
rect 103200 39448 104000 39568
rect 0 38768 800 38888
rect 0 38088 800 38208
rect 103200 38088 104000 38208
rect 0 37408 800 37528
rect 103200 37408 104000 37528
rect 103200 36728 104000 36848
rect 0 36048 800 36168
rect 103200 36048 104000 36168
rect 0 35368 800 35488
rect 103200 35368 104000 35488
rect 0 34688 800 34808
rect 103200 34688 104000 34808
rect 0 34008 800 34128
rect 103200 34008 104000 34128
rect 0 33328 800 33448
rect 103200 33328 104000 33448
rect 0 32648 800 32768
rect 103200 32648 104000 32768
rect 0 31968 800 32088
rect 103200 31968 104000 32088
rect 0 31288 800 31408
rect 103200 31288 104000 31408
rect 0 30608 800 30728
rect 103200 30608 104000 30728
rect 0 29928 800 30048
rect 103200 29928 104000 30048
rect 0 29248 800 29368
rect 103200 29248 104000 29368
rect 0 28568 800 28688
rect 103200 28568 104000 28688
rect 0 27888 800 28008
rect 103200 27888 104000 28008
rect 0 27208 800 27328
rect 103200 27208 104000 27328
rect 0 26528 800 26648
rect 103200 26528 104000 26648
rect 0 25848 800 25968
rect 103200 25848 104000 25968
rect 0 25168 800 25288
rect 103200 25168 104000 25288
rect 0 24488 800 24608
rect 103200 24488 104000 24608
rect 0 23808 800 23928
rect 103200 23808 104000 23928
rect 0 23128 800 23248
rect 103200 23128 104000 23248
rect 0 22448 800 22568
rect 103200 22448 104000 22568
rect 0 21768 800 21888
rect 103200 21768 104000 21888
rect 0 21088 800 21208
rect 103200 21088 104000 21208
rect 0 20408 800 20528
rect 103200 20408 104000 20528
rect 0 19728 800 19848
rect 0 19048 800 19168
rect 103200 19048 104000 19168
rect 103200 18368 104000 18488
rect 0 17688 800 17808
rect 103200 17688 104000 17808
rect 0 17008 800 17128
rect 103200 17008 104000 17128
rect 0 16328 800 16448
rect 103200 16328 104000 16448
rect 0 15648 800 15768
rect 103200 15648 104000 15768
rect 0 14968 800 15088
rect 103200 14968 104000 15088
rect 0 14288 800 14408
rect 103200 14288 104000 14408
rect 0 13608 800 13728
rect 103200 13608 104000 13728
rect 0 12928 800 13048
rect 103200 12928 104000 13048
rect 0 12248 800 12368
rect 103200 12248 104000 12368
rect 0 11568 800 11688
rect 103200 11568 104000 11688
rect 0 10888 800 11008
rect 103200 10888 104000 11008
rect 0 10208 800 10328
rect 103200 10208 104000 10328
rect 0 9528 800 9648
rect 103200 9528 104000 9648
rect 0 8848 800 8968
rect 103200 8848 104000 8968
rect 0 8168 800 8288
rect 103200 8168 104000 8288
rect 0 7488 800 7608
rect 103200 7488 104000 7608
rect 0 6808 800 6928
rect 103200 6808 104000 6928
rect 0 6128 800 6248
rect 103200 6128 104000 6248
rect 0 5448 800 5568
rect 103200 5448 104000 5568
rect 0 4768 800 4888
rect 103200 4768 104000 4888
rect 0 4088 800 4208
rect 103200 4088 104000 4208
rect 0 3408 800 3528
rect 103200 3408 104000 3528
rect 0 2728 800 2848
rect 103200 2728 104000 2848
rect 0 2048 800 2168
rect 103200 2048 104000 2168
rect 0 1368 800 1488
rect 0 688 800 808
rect 103200 688 104000 808
rect 103200 8 104000 128
<< obsm3 >>
rect 880 103288 103120 103461
rect 800 102888 103200 103288
rect 880 102608 103120 102888
rect 800 102208 103200 102608
rect 880 101928 103120 102208
rect 800 101528 103200 101928
rect 880 101248 103120 101528
rect 800 100848 103200 101248
rect 880 100568 103120 100848
rect 800 100168 103200 100568
rect 880 99888 103120 100168
rect 800 99488 103200 99888
rect 880 99208 103120 99488
rect 800 98808 103200 99208
rect 880 98528 103120 98808
rect 800 98128 103200 98528
rect 880 97848 103120 98128
rect 800 97448 103200 97848
rect 880 97168 103120 97448
rect 800 96768 103200 97168
rect 880 96488 103120 96768
rect 800 96088 103200 96488
rect 880 95808 103120 96088
rect 800 95408 103200 95808
rect 880 95128 103120 95408
rect 800 94728 103200 95128
rect 880 94448 103200 94728
rect 800 94048 103200 94448
rect 880 93768 103120 94048
rect 800 93368 103200 93768
rect 880 93088 103120 93368
rect 800 92688 103200 93088
rect 800 92408 103120 92688
rect 800 92008 103200 92408
rect 880 91728 103120 92008
rect 800 91328 103200 91728
rect 880 91048 103120 91328
rect 800 90648 103200 91048
rect 880 90368 103120 90648
rect 800 89968 103200 90368
rect 880 89688 103120 89968
rect 800 89288 103200 89688
rect 880 89008 103120 89288
rect 800 88608 103200 89008
rect 880 88328 103120 88608
rect 800 87928 103200 88328
rect 880 87648 103120 87928
rect 800 87248 103200 87648
rect 880 86968 103120 87248
rect 800 86568 103200 86968
rect 880 86288 103120 86568
rect 800 85888 103200 86288
rect 880 85608 103120 85888
rect 800 85208 103200 85608
rect 880 84928 103120 85208
rect 800 84528 103200 84928
rect 880 84248 103120 84528
rect 800 83848 103200 84248
rect 880 83568 103120 83848
rect 800 83168 103200 83568
rect 880 82888 103120 83168
rect 800 82488 103200 82888
rect 880 82208 103120 82488
rect 800 81808 103200 82208
rect 880 81528 103120 81808
rect 800 81128 103200 81528
rect 880 80848 103120 81128
rect 800 80448 103200 80848
rect 880 80168 103120 80448
rect 800 79768 103200 80168
rect 880 79488 103120 79768
rect 800 79088 103200 79488
rect 880 78808 103120 79088
rect 800 78408 103200 78808
rect 880 78128 103120 78408
rect 800 77728 103200 78128
rect 880 77448 103120 77728
rect 800 77048 103200 77448
rect 880 76768 103120 77048
rect 800 76368 103200 76768
rect 880 76088 103120 76368
rect 800 75688 103200 76088
rect 880 75408 103200 75688
rect 800 75008 103200 75408
rect 880 74728 103120 75008
rect 800 74328 103200 74728
rect 800 74048 103120 74328
rect 800 73648 103200 74048
rect 880 73368 103120 73648
rect 800 72968 103200 73368
rect 880 72688 103120 72968
rect 800 72288 103200 72688
rect 880 72008 103120 72288
rect 800 71608 103200 72008
rect 880 71328 103120 71608
rect 800 70928 103200 71328
rect 880 70648 103120 70928
rect 800 70248 103200 70648
rect 880 69968 103120 70248
rect 800 69568 103200 69968
rect 880 69288 103120 69568
rect 800 68888 103200 69288
rect 880 68608 103120 68888
rect 800 68208 103200 68608
rect 880 67928 103120 68208
rect 800 67528 103200 67928
rect 880 67248 103120 67528
rect 800 66848 103200 67248
rect 880 66568 103120 66848
rect 800 66168 103200 66568
rect 880 65888 103120 66168
rect 800 65488 103200 65888
rect 880 65208 103120 65488
rect 800 64808 103200 65208
rect 880 64528 103120 64808
rect 800 64128 103200 64528
rect 880 63848 103120 64128
rect 800 63448 103200 63848
rect 880 63168 103120 63448
rect 800 62768 103200 63168
rect 880 62488 103120 62768
rect 800 62088 103200 62488
rect 880 61808 103120 62088
rect 800 61408 103200 61808
rect 880 61128 103120 61408
rect 800 60728 103200 61128
rect 880 60448 103120 60728
rect 800 60048 103200 60448
rect 880 59768 103120 60048
rect 800 59368 103200 59768
rect 880 59088 103120 59368
rect 800 58688 103200 59088
rect 880 58408 103120 58688
rect 800 58008 103200 58408
rect 880 57728 103120 58008
rect 800 57328 103200 57728
rect 880 57048 103200 57328
rect 800 56648 103200 57048
rect 880 56368 103120 56648
rect 800 55968 103200 56368
rect 800 55688 103120 55968
rect 800 55288 103200 55688
rect 880 55008 103120 55288
rect 800 54608 103200 55008
rect 880 54328 103120 54608
rect 800 53928 103200 54328
rect 880 53648 103120 53928
rect 800 53248 103200 53648
rect 880 52968 103120 53248
rect 800 52568 103200 52968
rect 880 52288 103120 52568
rect 800 51888 103200 52288
rect 880 51608 103120 51888
rect 800 51208 103200 51608
rect 880 50928 103120 51208
rect 800 50528 103200 50928
rect 880 50248 103120 50528
rect 800 49848 103200 50248
rect 880 49568 103120 49848
rect 800 49168 103200 49568
rect 880 48888 103120 49168
rect 800 48488 103200 48888
rect 880 48208 103120 48488
rect 800 47808 103200 48208
rect 880 47528 103120 47808
rect 800 47128 103200 47528
rect 880 46848 103120 47128
rect 800 46448 103200 46848
rect 880 46168 103120 46448
rect 800 45768 103200 46168
rect 880 45488 103120 45768
rect 800 45088 103200 45488
rect 880 44808 103120 45088
rect 800 44408 103200 44808
rect 880 44128 103120 44408
rect 800 43728 103200 44128
rect 880 43448 103120 43728
rect 800 43048 103200 43448
rect 880 42768 103120 43048
rect 800 42368 103200 42768
rect 880 42088 103120 42368
rect 800 41688 103200 42088
rect 880 41408 103120 41688
rect 800 41008 103200 41408
rect 880 40728 103120 41008
rect 800 40328 103200 40728
rect 880 40048 103120 40328
rect 800 39648 103200 40048
rect 880 39368 103120 39648
rect 800 38968 103200 39368
rect 880 38688 103200 38968
rect 800 38288 103200 38688
rect 880 38008 103120 38288
rect 800 37608 103200 38008
rect 880 37328 103120 37608
rect 800 36928 103200 37328
rect 800 36648 103120 36928
rect 800 36248 103200 36648
rect 880 35968 103120 36248
rect 800 35568 103200 35968
rect 880 35288 103120 35568
rect 800 34888 103200 35288
rect 880 34608 103120 34888
rect 800 34208 103200 34608
rect 880 33928 103120 34208
rect 800 33528 103200 33928
rect 880 33248 103120 33528
rect 800 32848 103200 33248
rect 880 32568 103120 32848
rect 800 32168 103200 32568
rect 880 31888 103120 32168
rect 800 31488 103200 31888
rect 880 31208 103120 31488
rect 800 30808 103200 31208
rect 880 30528 103120 30808
rect 800 30128 103200 30528
rect 880 29848 103120 30128
rect 800 29448 103200 29848
rect 880 29168 103120 29448
rect 800 28768 103200 29168
rect 880 28488 103120 28768
rect 800 28088 103200 28488
rect 880 27808 103120 28088
rect 800 27408 103200 27808
rect 880 27128 103120 27408
rect 800 26728 103200 27128
rect 880 26448 103120 26728
rect 800 26048 103200 26448
rect 880 25768 103120 26048
rect 800 25368 103200 25768
rect 880 25088 103120 25368
rect 800 24688 103200 25088
rect 880 24408 103120 24688
rect 800 24008 103200 24408
rect 880 23728 103120 24008
rect 800 23328 103200 23728
rect 880 23048 103120 23328
rect 800 22648 103200 23048
rect 880 22368 103120 22648
rect 800 21968 103200 22368
rect 880 21688 103120 21968
rect 800 21288 103200 21688
rect 880 21008 103120 21288
rect 800 20608 103200 21008
rect 880 20328 103120 20608
rect 800 19928 103200 20328
rect 880 19648 103200 19928
rect 800 19248 103200 19648
rect 880 18968 103120 19248
rect 800 18568 103200 18968
rect 800 18288 103120 18568
rect 800 17888 103200 18288
rect 880 17608 103120 17888
rect 800 17208 103200 17608
rect 880 16928 103120 17208
rect 800 16528 103200 16928
rect 880 16248 103120 16528
rect 800 15848 103200 16248
rect 880 15568 103120 15848
rect 800 15168 103200 15568
rect 880 14888 103120 15168
rect 800 14488 103200 14888
rect 880 14208 103120 14488
rect 800 13808 103200 14208
rect 880 13528 103120 13808
rect 800 13128 103200 13528
rect 880 12848 103120 13128
rect 800 12448 103200 12848
rect 880 12168 103120 12448
rect 800 11768 103200 12168
rect 880 11488 103120 11768
rect 800 11088 103200 11488
rect 880 10808 103120 11088
rect 800 10408 103200 10808
rect 880 10128 103120 10408
rect 800 9728 103200 10128
rect 880 9448 103120 9728
rect 800 9048 103200 9448
rect 880 8768 103120 9048
rect 800 8368 103200 8768
rect 880 8088 103120 8368
rect 800 7688 103200 8088
rect 880 7408 103120 7688
rect 800 7008 103200 7408
rect 880 6728 103120 7008
rect 800 6328 103200 6728
rect 880 6048 103120 6328
rect 800 5648 103200 6048
rect 880 5368 103120 5648
rect 800 4968 103200 5368
rect 880 4688 103120 4968
rect 800 4288 103200 4688
rect 880 4008 103120 4288
rect 800 3608 103200 4008
rect 880 3328 103120 3608
rect 800 2928 103200 3328
rect 880 2648 103120 2928
rect 800 2248 103200 2648
rect 880 1968 103120 2248
rect 800 1568 103200 1968
rect 880 1288 103200 1568
rect 800 888 103200 1288
rect 880 608 103120 888
rect 800 208 103200 608
rect 800 35 103120 208
<< labels >>
rlabel metal2 s 4868 2128 5188 101776 6 VGND
port 1 nsew ground bidirectional
rlabel metal2 s 35588 2128 35908 101776 6 VGND
port 1 nsew ground bidirectional
rlabel metal2 s 66308 2128 66628 101776 6 VGND
port 1 nsew ground bidirectional
rlabel metal2 s 97028 2128 97348 101776 6 VGND
port 1 nsew ground bidirectional
rlabel metal2 s 4208 2128 4528 101776 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 34928 2128 35248 101776 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 65648 2128 65968 101776 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 96368 2128 96688 101776 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 99194 0 99250 800 6 io_in[0]
port 3 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 103200 44888 104000 45008 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 io_in[12]
port 6 nsew signal input
rlabel metal2 s 35438 103200 35494 104000 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 103200 67328 104000 67448 6 io_in[14]
port 8 nsew signal input
rlabel metal2 s 30286 103200 30342 104000 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 103200 99288 104000 99408 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_in[18]
port 12 nsew signal input
rlabel metal2 s 38658 103200 38714 104000 6 io_in[19]
port 13 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_in[1]
port 14 nsew signal input
rlabel metal2 s 27066 103200 27122 104000 6 io_in[20]
port 15 nsew signal input
rlabel metal2 s 32218 103200 32274 104000 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 103200 76848 104000 76968 6 io_in[24]
port 19 nsew signal input
rlabel metal2 s 4526 103200 4582 104000 6 io_in[25]
port 20 nsew signal input
rlabel metal2 s 65706 103200 65762 104000 6 io_in[26]
port 21 nsew signal input
rlabel metal2 s 28998 103200 29054 104000 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_in[28]
port 23 nsew signal input
rlabel metal2 s 47674 103200 47730 104000 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 io_in[2]
port 25 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_in[31]
port 27 nsew signal input
rlabel metal2 s 70858 103200 70914 104000 6 io_in[32]
port 28 nsew signal input
rlabel metal2 s 61198 103200 61254 104000 6 io_in[33]
port 29 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 io_in[34]
port 30 nsew signal input
rlabel metal3 s 103200 68008 104000 68128 6 io_in[35]
port 31 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 io_in[36]
port 32 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 io_in[37]
port 33 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 io_in[3]
port 34 nsew signal input
rlabel metal2 s 98550 103200 98606 104000 6 io_in[4]
port 35 nsew signal input
rlabel metal3 s 103200 10888 104000 11008 6 io_in[5]
port 36 nsew signal input
rlabel metal3 s 103200 60528 104000 60648 6 io_in[6]
port 37 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 io_in[7]
port 38 nsew signal input
rlabel metal2 s 50250 103200 50306 104000 6 io_in[8]
port 39 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 io_in[9]
port 40 nsew signal input
rlabel metal3 s 103200 35368 104000 35488 6 io_oeb[0]
port 41 nsew signal output
rlabel metal3 s 103200 33328 104000 33448 6 io_oeb[10]
port 42 nsew signal output
rlabel metal2 s 62486 103200 62542 104000 6 io_oeb[11]
port 43 nsew signal output
rlabel metal2 s 36726 103200 36782 104000 6 io_oeb[12]
port 44 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 io_oeb[13]
port 45 nsew signal output
rlabel metal2 s 18694 103200 18750 104000 6 io_oeb[14]
port 46 nsew signal output
rlabel metal3 s 103200 36048 104000 36168 6 io_oeb[15]
port 47 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 io_oeb[16]
port 48 nsew signal output
rlabel metal2 s 1306 103200 1362 104000 6 io_oeb[17]
port 49 nsew signal output
rlabel metal2 s 3238 103200 3294 104000 6 io_oeb[18]
port 50 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_oeb[19]
port 51 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 io_oeb[1]
port 52 nsew signal output
rlabel metal2 s 19338 103200 19394 104000 6 io_oeb[20]
port 53 nsew signal output
rlabel metal2 s 71502 103200 71558 104000 6 io_oeb[21]
port 54 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 io_oeb[22]
port 55 nsew signal output
rlabel metal3 s 103200 41488 104000 41608 6 io_oeb[23]
port 56 nsew signal output
rlabel metal3 s 103200 102688 104000 102808 6 io_oeb[24]
port 57 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 io_oeb[25]
port 58 nsew signal output
rlabel metal2 s 12898 103200 12954 104000 6 io_oeb[26]
port 59 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_oeb[27]
port 60 nsew signal output
rlabel metal2 s 63774 103200 63830 104000 6 io_oeb[28]
port 61 nsew signal output
rlabel metal3 s 103200 76168 104000 76288 6 io_oeb[29]
port 62 nsew signal output
rlabel metal3 s 103200 89088 104000 89208 6 io_oeb[2]
port 63 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 io_oeb[30]
port 64 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 io_oeb[31]
port 65 nsew signal output
rlabel metal2 s 14186 103200 14242 104000 6 io_oeb[32]
port 66 nsew signal output
rlabel metal2 s 5170 103200 5226 104000 6 io_oeb[33]
port 67 nsew signal output
rlabel metal2 s 19982 103200 20038 104000 6 io_oeb[34]
port 68 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 io_oeb[35]
port 69 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 io_oeb[36]
port 70 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 io_oeb[37]
port 71 nsew signal output
rlabel metal2 s 79874 103200 79930 104000 6 io_oeb[3]
port 72 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 io_oeb[4]
port 73 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_oeb[5]
port 74 nsew signal output
rlabel metal2 s 74722 103200 74778 104000 6 io_oeb[6]
port 75 nsew signal output
rlabel metal2 s 100482 103200 100538 104000 6 io_oeb[7]
port 76 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 io_oeb[8]
port 77 nsew signal output
rlabel metal2 s 11610 103200 11666 104000 6 io_oeb[9]
port 78 nsew signal output
rlabel metal2 s 18 103200 74 104000 6 io_out[0]
port 79 nsew signal output
rlabel metal2 s 97906 103200 97962 104000 6 io_out[10]
port 80 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_out[11]
port 81 nsew signal output
rlabel metal3 s 103200 96568 104000 96688 6 io_out[12]
port 82 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 io_out[13]
port 83 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 io_out[14]
port 84 nsew signal output
rlabel metal3 s 103200 80248 104000 80368 6 io_out[15]
port 85 nsew signal output
rlabel metal3 s 103200 22448 104000 22568 6 io_out[16]
port 86 nsew signal output
rlabel metal3 s 103200 66648 104000 66768 6 io_out[17]
port 87 nsew signal output
rlabel metal3 s 103200 92488 104000 92608 6 io_out[18]
port 88 nsew signal output
rlabel metal3 s 103200 80928 104000 81048 6 io_out[19]
port 89 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 io_out[1]
port 90 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 io_out[20]
port 91 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 io_out[21]
port 92 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 io_out[22]
port 93 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 io_out[23]
port 94 nsew signal output
rlabel metal3 s 103200 9528 104000 9648 6 io_out[24]
port 95 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 io_out[25]
port 96 nsew signal output
rlabel metal2 s 21270 103200 21326 104000 6 io_out[26]
port 97 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 io_out[27]
port 98 nsew signal output
rlabel metal3 s 103200 56448 104000 56568 6 io_out[28]
port 99 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 io_out[29]
port 100 nsew signal output
rlabel metal2 s 99838 103200 99894 104000 6 io_out[2]
port 101 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 io_out[30]
port 102 nsew signal output
rlabel metal3 s 103200 91128 104000 91248 6 io_out[31]
port 103 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 io_out[32]
port 104 nsew signal output
rlabel metal3 s 103200 78208 104000 78328 6 io_out[33]
port 105 nsew signal output
rlabel metal2 s 103058 103200 103114 104000 6 io_out[34]
port 106 nsew signal output
rlabel metal3 s 103200 69368 104000 69488 6 io_out[35]
port 107 nsew signal output
rlabel metal2 s 20626 103200 20682 104000 6 io_out[36]
port 108 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 io_out[37]
port 109 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 io_out[3]
port 110 nsew signal output
rlabel metal3 s 103200 8168 104000 8288 6 io_out[4]
port 111 nsew signal output
rlabel metal3 s 103200 63928 104000 64048 6 io_out[5]
port 112 nsew signal output
rlabel metal2 s 52826 103200 52882 104000 6 io_out[6]
port 113 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_out[7]
port 114 nsew signal output
rlabel metal2 s 43166 103200 43222 104000 6 io_out[8]
port 115 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 io_out[9]
port 116 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 irq[0]
port 117 nsew signal output
rlabel metal3 s 103200 40808 104000 40928 6 irq[1]
port 118 nsew signal output
rlabel metal2 s 82450 103200 82506 104000 6 irq[2]
port 119 nsew signal output
rlabel metal3 s 103200 51688 104000 51808 6 la_data_in[0]
port 120 nsew signal input
rlabel metal3 s 103200 27888 104000 28008 6 la_data_in[100]
port 121 nsew signal input
rlabel metal2 s 46386 103200 46442 104000 6 la_data_in[101]
port 122 nsew signal input
rlabel metal2 s 17406 103200 17462 104000 6 la_data_in[102]
port 123 nsew signal input
rlabel metal3 s 103200 95208 104000 95328 6 la_data_in[103]
port 124 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_data_in[104]
port 125 nsew signal input
rlabel metal3 s 103200 64608 104000 64728 6 la_data_in[105]
port 126 nsew signal input
rlabel metal3 s 103200 8848 104000 8968 6 la_data_in[106]
port 127 nsew signal input
rlabel metal2 s 56690 103200 56746 104000 6 la_data_in[107]
port 128 nsew signal input
rlabel metal3 s 103200 25848 104000 25968 6 la_data_in[108]
port 129 nsew signal input
rlabel metal2 s 74078 103200 74134 104000 6 la_data_in[109]
port 130 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 la_data_in[10]
port 131 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[110]
port 132 nsew signal input
rlabel metal3 s 103200 65288 104000 65408 6 la_data_in[111]
port 133 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 la_data_in[112]
port 134 nsew signal input
rlabel metal3 s 103200 14288 104000 14408 6 la_data_in[113]
port 135 nsew signal input
rlabel metal2 s 76654 103200 76710 104000 6 la_data_in[114]
port 136 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_data_in[115]
port 137 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[116]
port 138 nsew signal input
rlabel metal2 s 41878 103200 41934 104000 6 la_data_in[117]
port 139 nsew signal input
rlabel metal2 s 83738 103200 83794 104000 6 la_data_in[118]
port 140 nsew signal input
rlabel metal3 s 103200 61888 104000 62008 6 la_data_in[119]
port 141 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 la_data_in[11]
port 142 nsew signal input
rlabel metal2 s 70214 103200 70270 104000 6 la_data_in[120]
port 143 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[121]
port 144 nsew signal input
rlabel metal2 s 5814 103200 5870 104000 6 la_data_in[122]
port 145 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[123]
port 146 nsew signal input
rlabel metal2 s 10322 103200 10378 104000 6 la_data_in[124]
port 147 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 la_data_in[125]
port 148 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[126]
port 149 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_data_in[127]
port 150 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 la_data_in[12]
port 151 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[13]
port 152 nsew signal input
rlabel metal3 s 103200 74128 104000 74248 6 la_data_in[14]
port 153 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 la_data_in[15]
port 154 nsew signal input
rlabel metal3 s 103200 42848 104000 42968 6 la_data_in[16]
port 155 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 la_data_in[17]
port 156 nsew signal input
rlabel metal3 s 103200 87048 104000 87168 6 la_data_in[18]
port 157 nsew signal input
rlabel metal2 s 79230 103200 79286 104000 6 la_data_in[19]
port 158 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_data_in[1]
port 159 nsew signal input
rlabel metal2 s 2594 103200 2650 104000 6 la_data_in[20]
port 160 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_data_in[21]
port 161 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[22]
port 162 nsew signal input
rlabel metal3 s 103200 53728 104000 53848 6 la_data_in[23]
port 163 nsew signal input
rlabel metal3 s 103200 18368 104000 18488 6 la_data_in[24]
port 164 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 la_data_in[25]
port 165 nsew signal input
rlabel metal3 s 103200 82968 104000 83088 6 la_data_in[26]
port 166 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 la_data_in[27]
port 167 nsew signal input
rlabel metal3 s 103200 61208 104000 61328 6 la_data_in[28]
port 168 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[29]
port 169 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[2]
port 170 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[30]
port 171 nsew signal input
rlabel metal2 s 38014 103200 38070 104000 6 la_data_in[31]
port 172 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[32]
port 173 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[33]
port 174 nsew signal input
rlabel metal2 s 48318 103200 48374 104000 6 la_data_in[34]
port 175 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 la_data_in[35]
port 176 nsew signal input
rlabel metal2 s 81806 103200 81862 104000 6 la_data_in[36]
port 177 nsew signal input
rlabel metal2 s 101126 103200 101182 104000 6 la_data_in[37]
port 178 nsew signal input
rlabel metal3 s 103200 44208 104000 44328 6 la_data_in[38]
port 179 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 la_data_in[39]
port 180 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_data_in[3]
port 181 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_data_in[40]
port 182 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[41]
port 183 nsew signal input
rlabel metal3 s 103200 46248 104000 46368 6 la_data_in[42]
port 184 nsew signal input
rlabel metal3 s 103200 79568 104000 79688 6 la_data_in[43]
port 185 nsew signal input
rlabel metal2 s 34794 103200 34850 104000 6 la_data_in[44]
port 186 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_data_in[45]
port 187 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 la_data_in[46]
port 188 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[47]
port 189 nsew signal input
rlabel metal2 s 73434 103200 73490 104000 6 la_data_in[48]
port 190 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_data_in[49]
port 191 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[4]
port 192 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 la_data_in[50]
port 193 nsew signal input
rlabel metal2 s 1950 103200 2006 104000 6 la_data_in[51]
port 194 nsew signal input
rlabel metal2 s 99194 103200 99250 104000 6 la_data_in[52]
port 195 nsew signal input
rlabel metal3 s 103200 17688 104000 17808 6 la_data_in[53]
port 196 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_data_in[54]
port 197 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[55]
port 198 nsew signal input
rlabel metal2 s 662 0 718 800 6 la_data_in[56]
port 199 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[57]
port 200 nsew signal input
rlabel metal2 s 86314 103200 86370 104000 6 la_data_in[58]
port 201 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[59]
port 202 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 la_data_in[5]
port 203 nsew signal input
rlabel metal2 s 9034 103200 9090 104000 6 la_data_in[60]
port 204 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_data_in[61]
port 205 nsew signal input
rlabel metal3 s 103200 23808 104000 23928 6 la_data_in[62]
port 206 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 la_data_in[63]
port 207 nsew signal input
rlabel metal3 s 103200 97928 104000 98048 6 la_data_in[64]
port 208 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[65]
port 209 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 la_data_in[66]
port 210 nsew signal input
rlabel metal2 s 43810 103200 43866 104000 6 la_data_in[67]
port 211 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 la_data_in[68]
port 212 nsew signal input
rlabel metal3 s 103200 74808 104000 74928 6 la_data_in[69]
port 213 nsew signal input
rlabel metal3 s 103200 40128 104000 40248 6 la_data_in[6]
port 214 nsew signal input
rlabel metal3 s 103200 24488 104000 24608 6 la_data_in[70]
port 215 nsew signal input
rlabel metal3 s 103200 17008 104000 17128 6 la_data_in[71]
port 216 nsew signal input
rlabel metal2 s 26422 103200 26478 104000 6 la_data_in[72]
port 217 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_data_in[73]
port 218 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[74]
port 219 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[75]
port 220 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[76]
port 221 nsew signal input
rlabel metal3 s 103200 65968 104000 66088 6 la_data_in[77]
port 222 nsew signal input
rlabel metal3 s 103200 82288 104000 82408 6 la_data_in[78]
port 223 nsew signal input
rlabel metal3 s 103200 27208 104000 27328 6 la_data_in[79]
port 224 nsew signal input
rlabel metal3 s 103200 30608 104000 30728 6 la_data_in[7]
port 225 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[80]
port 226 nsew signal input
rlabel metal3 s 103200 31288 104000 31408 6 la_data_in[81]
port 227 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 la_data_in[82]
port 228 nsew signal input
rlabel metal2 s 86958 103200 87014 104000 6 la_data_in[83]
port 229 nsew signal input
rlabel metal3 s 0 688 800 808 6 la_data_in[84]
port 230 nsew signal input
rlabel metal2 s 41234 103200 41290 104000 6 la_data_in[85]
port 231 nsew signal input
rlabel metal3 s 103200 72768 104000 72888 6 la_data_in[86]
port 232 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 la_data_in[87]
port 233 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 la_data_in[88]
port 234 nsew signal input
rlabel metal2 s 36082 103200 36138 104000 6 la_data_in[89]
port 235 nsew signal input
rlabel metal2 s 25134 103200 25190 104000 6 la_data_in[8]
port 236 nsew signal input
rlabel metal2 s 60554 103200 60610 104000 6 la_data_in[90]
port 237 nsew signal input
rlabel metal2 s 3882 103200 3938 104000 6 la_data_in[91]
port 238 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[92]
port 239 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[93]
port 240 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[94]
port 241 nsew signal input
rlabel metal3 s 103200 6808 104000 6928 6 la_data_in[95]
port 242 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_data_in[96]
port 243 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 la_data_in[97]
port 244 nsew signal input
rlabel metal3 s 103200 47608 104000 47728 6 la_data_in[98]
port 245 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_data_in[99]
port 246 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 la_data_in[9]
port 247 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 la_data_out[0]
port 248 nsew signal output
rlabel metal2 s 96618 103200 96674 104000 6 la_data_out[100]
port 249 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 la_data_out[101]
port 250 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 la_data_out[102]
port 251 nsew signal output
rlabel metal3 s 103200 36728 104000 36848 6 la_data_out[103]
port 252 nsew signal output
rlabel metal3 s 103200 55088 104000 55208 6 la_data_out[104]
port 253 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 la_data_out[105]
port 254 nsew signal output
rlabel metal2 s 23846 103200 23902 104000 6 la_data_out[106]
port 255 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[107]
port 256 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 la_data_out[108]
port 257 nsew signal output
rlabel metal2 s 54114 103200 54170 104000 6 la_data_out[109]
port 258 nsew signal output
rlabel metal2 s 63130 103200 63186 104000 6 la_data_out[10]
port 259 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 la_data_out[110]
port 260 nsew signal output
rlabel metal2 s 76010 103200 76066 104000 6 la_data_out[111]
port 261 nsew signal output
rlabel metal2 s 94042 103200 94098 104000 6 la_data_out[112]
port 262 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 la_data_out[113]
port 263 nsew signal output
rlabel metal2 s 44454 103200 44510 104000 6 la_data_out[114]
port 264 nsew signal output
rlabel metal3 s 103200 90448 104000 90568 6 la_data_out[115]
port 265 nsew signal output
rlabel metal3 s 103200 21768 104000 21888 6 la_data_out[116]
port 266 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 la_data_out[117]
port 267 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_data_out[118]
port 268 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 la_data_out[119]
port 269 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[11]
port 270 nsew signal output
rlabel metal3 s 103200 688 104000 808 6 la_data_out[120]
port 271 nsew signal output
rlabel metal2 s 18050 103200 18106 104000 6 la_data_out[121]
port 272 nsew signal output
rlabel metal2 s 95974 103200 96030 104000 6 la_data_out[122]
port 273 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 la_data_out[123]
port 274 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 la_data_out[124]
port 275 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[125]
port 276 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[126]
port 277 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 la_data_out[127]
port 278 nsew signal output
rlabel metal3 s 103200 91808 104000 91928 6 la_data_out[12]
port 279 nsew signal output
rlabel metal3 s 103200 45568 104000 45688 6 la_data_out[13]
port 280 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 la_data_out[14]
port 281 nsew signal output
rlabel metal3 s 103200 50328 104000 50448 6 la_data_out[15]
port 282 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[16]
port 283 nsew signal output
rlabel metal2 s 9678 103200 9734 104000 6 la_data_out[17]
port 284 nsew signal output
rlabel metal3 s 103200 15648 104000 15768 6 la_data_out[18]
port 285 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 la_data_out[19]
port 286 nsew signal output
rlabel metal2 s 8390 103200 8446 104000 6 la_data_out[1]
port 287 nsew signal output
rlabel metal3 s 103200 100648 104000 100768 6 la_data_out[20]
port 288 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 la_data_out[21]
port 289 nsew signal output
rlabel metal2 s 68282 103200 68338 104000 6 la_data_out[22]
port 290 nsew signal output
rlabel metal3 s 103200 37408 104000 37528 6 la_data_out[23]
port 291 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 la_data_out[24]
port 292 nsew signal output
rlabel metal2 s 57978 103200 58034 104000 6 la_data_out[25]
port 293 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 la_data_out[26]
port 294 nsew signal output
rlabel metal3 s 103200 46928 104000 47048 6 la_data_out[27]
port 295 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 la_data_out[28]
port 296 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 la_data_out[29]
port 297 nsew signal output
rlabel metal3 s 103200 12928 104000 13048 6 la_data_out[2]
port 298 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[30]
port 299 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out[31]
port 300 nsew signal output
rlabel metal2 s 22558 103200 22614 104000 6 la_data_out[32]
port 301 nsew signal output
rlabel metal2 s 59266 103200 59322 104000 6 la_data_out[33]
port 302 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[34]
port 303 nsew signal output
rlabel metal2 s 91466 103200 91522 104000 6 la_data_out[35]
port 304 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 la_data_out[36]
port 305 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 la_data_out[37]
port 306 nsew signal output
rlabel metal2 s 83094 103200 83150 104000 6 la_data_out[38]
port 307 nsew signal output
rlabel metal3 s 103200 26528 104000 26648 6 la_data_out[39]
port 308 nsew signal output
rlabel metal2 s 39946 103200 40002 104000 6 la_data_out[3]
port 309 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 la_data_out[40]
port 310 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[41]
port 311 nsew signal output
rlabel metal2 s 32862 103200 32918 104000 6 la_data_out[42]
port 312 nsew signal output
rlabel metal2 s 29642 103200 29698 104000 6 la_data_out[43]
port 313 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[44]
port 314 nsew signal output
rlabel metal3 s 103200 8 104000 128 6 la_data_out[45]
port 315 nsew signal output
rlabel metal2 s 102414 103200 102470 104000 6 la_data_out[46]
port 316 nsew signal output
rlabel metal2 s 37370 103200 37426 104000 6 la_data_out[47]
port 317 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 la_data_out[48]
port 318 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 la_data_out[49]
port 319 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 la_data_out[4]
port 320 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 la_data_out[50]
port 321 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[51]
port 322 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 la_data_out[52]
port 323 nsew signal output
rlabel metal3 s 103200 51008 104000 51128 6 la_data_out[53]
port 324 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 la_data_out[54]
port 325 nsew signal output
rlabel metal3 s 103200 48288 104000 48408 6 la_data_out[55]
port 326 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 la_data_out[56]
port 327 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[57]
port 328 nsew signal output
rlabel metal2 s 97262 103200 97318 104000 6 la_data_out[58]
port 329 nsew signal output
rlabel metal2 s 80518 103200 80574 104000 6 la_data_out[59]
port 330 nsew signal output
rlabel metal2 s 50894 103200 50950 104000 6 la_data_out[5]
port 331 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 la_data_out[60]
port 332 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[61]
port 333 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 la_data_out[62]
port 334 nsew signal output
rlabel metal3 s 103200 54408 104000 54528 6 la_data_out[63]
port 335 nsew signal output
rlabel metal3 s 103200 21088 104000 21208 6 la_data_out[64]
port 336 nsew signal output
rlabel metal3 s 103200 11568 104000 11688 6 la_data_out[65]
port 337 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[66]
port 338 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[67]
port 339 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[68]
port 340 nsew signal output
rlabel metal2 s 93398 103200 93454 104000 6 la_data_out[69]
port 341 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[6]
port 342 nsew signal output
rlabel metal2 s 40590 103200 40646 104000 6 la_data_out[70]
port 343 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 la_data_out[71]
port 344 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 la_data_out[72]
port 345 nsew signal output
rlabel metal2 s 52182 103200 52238 104000 6 la_data_out[73]
port 346 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 la_data_out[74]
port 347 nsew signal output
rlabel metal3 s 103200 7488 104000 7608 6 la_data_out[75]
port 348 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[76]
port 349 nsew signal output
rlabel metal3 s 103200 20408 104000 20528 6 la_data_out[77]
port 350 nsew signal output
rlabel metal3 s 103200 14968 104000 15088 6 la_data_out[78]
port 351 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[79]
port 352 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 la_data_out[7]
port 353 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 la_data_out[80]
port 354 nsew signal output
rlabel metal2 s 23202 103200 23258 104000 6 la_data_out[81]
port 355 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[82]
port 356 nsew signal output
rlabel metal2 s 16118 103200 16174 104000 6 la_data_out[83]
port 357 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[84]
port 358 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 la_data_out[85]
port 359 nsew signal output
rlabel metal3 s 103200 52368 104000 52488 6 la_data_out[86]
port 360 nsew signal output
rlabel metal2 s 57334 103200 57390 104000 6 la_data_out[87]
port 361 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[88]
port 362 nsew signal output
rlabel metal2 s 54758 103200 54814 104000 6 la_data_out[89]
port 363 nsew signal output
rlabel metal2 s 55402 103200 55458 104000 6 la_data_out[8]
port 364 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[90]
port 365 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[91]
port 366 nsew signal output
rlabel metal2 s 88246 103200 88302 104000 6 la_data_out[92]
port 367 nsew signal output
rlabel metal2 s 34150 103200 34206 104000 6 la_data_out[93]
port 368 nsew signal output
rlabel metal2 s 45098 103200 45154 104000 6 la_data_out[94]
port 369 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[95]
port 370 nsew signal output
rlabel metal2 s 10966 103200 11022 104000 6 la_data_out[96]
port 371 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la_data_out[97]
port 372 nsew signal output
rlabel metal2 s 85670 103200 85726 104000 6 la_data_out[98]
port 373 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[99]
port 374 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[9]
port 375 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 la_oenb[0]
port 376 nsew signal input
rlabel metal3 s 103200 102008 104000 102128 6 la_oenb[100]
port 377 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 la_oenb[101]
port 378 nsew signal input
rlabel metal2 s 87602 103200 87658 104000 6 la_oenb[102]
port 379 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_oenb[103]
port 380 nsew signal input
rlabel metal3 s 103200 59168 104000 59288 6 la_oenb[104]
port 381 nsew signal input
rlabel metal2 s 48962 103200 49018 104000 6 la_oenb[105]
port 382 nsew signal input
rlabel metal2 s 101770 103200 101826 104000 6 la_oenb[106]
port 383 nsew signal input
rlabel metal3 s 103200 57808 104000 57928 6 la_oenb[107]
port 384 nsew signal input
rlabel metal2 s 68926 103200 68982 104000 6 la_oenb[108]
port 385 nsew signal input
rlabel metal2 s 81162 103200 81218 104000 6 la_oenb[109]
port 386 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[10]
port 387 nsew signal input
rlabel metal3 s 103200 78888 104000 79008 6 la_oenb[110]
port 388 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[111]
port 389 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 la_oenb[112]
port 390 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_oenb[113]
port 391 nsew signal input
rlabel metal2 s 61842 103200 61898 104000 6 la_oenb[114]
port 392 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_oenb[115]
port 393 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[116]
port 394 nsew signal input
rlabel metal3 s 103200 98608 104000 98728 6 la_oenb[117]
port 395 nsew signal input
rlabel metal3 s 103200 39448 104000 39568 6 la_oenb[118]
port 396 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 la_oenb[119]
port 397 nsew signal input
rlabel metal3 s 103200 58488 104000 58608 6 la_oenb[11]
port 398 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[120]
port 399 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[121]
port 400 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 la_oenb[122]
port 401 nsew signal input
rlabel metal3 s 103200 85688 104000 85808 6 la_oenb[123]
port 402 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 la_oenb[124]
port 403 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 la_oenb[125]
port 404 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[126]
port 405 nsew signal input
rlabel metal3 s 103200 25168 104000 25288 6 la_oenb[127]
port 406 nsew signal input
rlabel metal3 s 103200 70728 104000 70848 6 la_oenb[12]
port 407 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_oenb[13]
port 408 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 la_oenb[14]
port 409 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[15]
port 410 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_oenb[16]
port 411 nsew signal input
rlabel metal3 s 103200 16328 104000 16448 6 la_oenb[17]
port 412 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 la_oenb[18]
port 413 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_oenb[19]
port 414 nsew signal input
rlabel metal3 s 103200 13608 104000 13728 6 la_oenb[1]
port 415 nsew signal input
rlabel metal3 s 103200 97248 104000 97368 6 la_oenb[20]
port 416 nsew signal input
rlabel metal3 s 103200 42168 104000 42288 6 la_oenb[21]
port 417 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 la_oenb[22]
port 418 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la_oenb[23]
port 419 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oenb[24]
port 420 nsew signal input
rlabel metal2 s 90822 103200 90878 104000 6 la_oenb[25]
port 421 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_oenb[26]
port 422 nsew signal input
rlabel metal3 s 103200 55768 104000 55888 6 la_oenb[27]
port 423 nsew signal input
rlabel metal2 s 103702 103200 103758 104000 6 la_oenb[28]
port 424 nsew signal input
rlabel metal2 s 92110 103200 92166 104000 6 la_oenb[29]
port 425 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_oenb[2]
port 426 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 la_oenb[30]
port 427 nsew signal input
rlabel metal2 s 30930 103200 30986 104000 6 la_oenb[31]
port 428 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[32]
port 429 nsew signal input
rlabel metal2 s 13542 103200 13598 104000 6 la_oenb[33]
port 430 nsew signal input
rlabel metal3 s 103200 31968 104000 32088 6 la_oenb[34]
port 431 nsew signal input
rlabel metal3 s 103200 59848 104000 59968 6 la_oenb[35]
port 432 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 la_oenb[36]
port 433 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oenb[37]
port 434 nsew signal input
rlabel metal3 s 103200 84328 104000 84448 6 la_oenb[38]
port 435 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_oenb[39]
port 436 nsew signal input
rlabel metal2 s 94686 103200 94742 104000 6 la_oenb[3]
port 437 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 la_oenb[40]
port 438 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[41]
port 439 nsew signal input
rlabel metal2 s 6458 103200 6514 104000 6 la_oenb[42]
port 440 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_oenb[43]
port 441 nsew signal input
rlabel metal3 s 103200 4768 104000 4888 6 la_oenb[44]
port 442 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_oenb[45]
port 443 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[46]
port 444 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[47]
port 445 nsew signal input
rlabel metal3 s 103200 29928 104000 30048 6 la_oenb[48]
port 446 nsew signal input
rlabel metal3 s 103200 85008 104000 85128 6 la_oenb[49]
port 447 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 la_oenb[4]
port 448 nsew signal input
rlabel metal2 s 49606 103200 49662 104000 6 la_oenb[50]
port 449 nsew signal input
rlabel metal2 s 33506 103200 33562 104000 6 la_oenb[51]
port 450 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 la_oenb[52]
port 451 nsew signal input
rlabel metal3 s 103200 95888 104000 96008 6 la_oenb[53]
port 452 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 la_oenb[54]
port 453 nsew signal input
rlabel metal2 s 27710 103200 27766 104000 6 la_oenb[55]
port 454 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 la_oenb[56]
port 455 nsew signal input
rlabel metal3 s 103200 83648 104000 83768 6 la_oenb[57]
port 456 nsew signal input
rlabel metal2 s 72790 103200 72846 104000 6 la_oenb[58]
port 457 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 la_oenb[59]
port 458 nsew signal input
rlabel metal2 s 84382 103200 84438 104000 6 la_oenb[5]
port 459 nsew signal input
rlabel metal2 s 89534 103200 89590 104000 6 la_oenb[60]
port 460 nsew signal input
rlabel metal2 s 90178 103200 90234 104000 6 la_oenb[61]
port 461 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[62]
port 462 nsew signal input
rlabel metal2 s 56046 103200 56102 104000 6 la_oenb[63]
port 463 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 la_oenb[64]
port 464 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la_oenb[65]
port 465 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[66]
port 466 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_oenb[67]
port 467 nsew signal input
rlabel metal3 s 103200 19048 104000 19168 6 la_oenb[68]
port 468 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 la_oenb[69]
port 469 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 la_oenb[6]
port 470 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 la_oenb[70]
port 471 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 la_oenb[71]
port 472 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_oenb[72]
port 473 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la_oenb[73]
port 474 nsew signal input
rlabel metal2 s 53470 103200 53526 104000 6 la_oenb[74]
port 475 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[75]
port 476 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[76]
port 477 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 la_oenb[77]
port 478 nsew signal input
rlabel metal3 s 103200 71408 104000 71528 6 la_oenb[78]
port 479 nsew signal input
rlabel metal3 s 103200 93848 104000 93968 6 la_oenb[79]
port 480 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_oenb[7]
port 481 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 la_oenb[80]
port 482 nsew signal input
rlabel metal3 s 103200 10208 104000 10328 6 la_oenb[81]
port 483 nsew signal input
rlabel metal3 s 103200 88408 104000 88528 6 la_oenb[82]
port 484 nsew signal input
rlabel metal2 s 39302 103200 39358 104000 6 la_oenb[83]
port 485 nsew signal input
rlabel metal3 s 103200 73448 104000 73568 6 la_oenb[84]
port 486 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[85]
port 487 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_oenb[86]
port 488 nsew signal input
rlabel metal3 s 103200 23128 104000 23248 6 la_oenb[87]
port 489 nsew signal input
rlabel metal2 s 31574 103200 31630 104000 6 la_oenb[88]
port 490 nsew signal input
rlabel metal3 s 103200 2048 104000 2168 6 la_oenb[89]
port 491 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 la_oenb[8]
port 492 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 la_oenb[90]
port 493 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 la_oenb[91]
port 494 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[92]
port 495 nsew signal input
rlabel metal3 s 103200 87728 104000 87848 6 la_oenb[93]
port 496 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_oenb[94]
port 497 nsew signal input
rlabel metal3 s 103200 3408 104000 3528 6 la_oenb[95]
port 498 nsew signal input
rlabel metal2 s 662 103200 718 104000 6 la_oenb[96]
port 499 nsew signal input
rlabel metal2 s 65062 103200 65118 104000 6 la_oenb[97]
port 500 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[98]
port 501 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 la_oenb[99]
port 502 nsew signal input
rlabel metal2 s 7746 103200 7802 104000 6 la_oenb[9]
port 503 nsew signal input
rlabel metal2 s 5528 2128 5848 101776 6 vccd1
port 504 nsew power bidirectional
rlabel metal2 s 36248 2128 36568 101776 6 vccd1
port 504 nsew power bidirectional
rlabel metal2 s 66968 2128 67288 101776 6 vccd1
port 504 nsew power bidirectional
rlabel metal2 s 97688 2128 98008 101776 6 vccd1
port 504 nsew power bidirectional
rlabel metal2 s 6188 2128 6508 101776 6 vssd1
port 505 nsew ground bidirectional
rlabel metal2 s 36908 2128 37228 101776 6 vssd1
port 505 nsew ground bidirectional
rlabel metal2 s 67628 2128 67948 101776 6 vssd1
port 505 nsew ground bidirectional
rlabel metal2 s 98348 2128 98668 101776 6 vssd1
port 505 nsew ground bidirectional
rlabel metal3 s 103200 29248 104000 29368 6 wb_clk_i
port 506 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 wb_rst_i
port 507 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wbs_ack_o
port 508 nsew signal output
rlabel metal2 s 45742 103200 45798 104000 6 wbs_adr_i[0]
port 509 nsew signal input
rlabel metal2 s 21914 103200 21970 104000 6 wbs_adr_i[10]
port 510 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 wbs_adr_i[11]
port 511 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[12]
port 512 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 wbs_adr_i[13]
port 513 nsew signal input
rlabel metal3 s 103200 93168 104000 93288 6 wbs_adr_i[14]
port 514 nsew signal input
rlabel metal3 s 103200 86368 104000 86488 6 wbs_adr_i[15]
port 515 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_adr_i[16]
port 516 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wbs_adr_i[17]
port 517 nsew signal input
rlabel metal3 s 103200 43528 104000 43648 6 wbs_adr_i[18]
port 518 nsew signal input
rlabel metal3 s 103200 2728 104000 2848 6 wbs_adr_i[19]
port 519 nsew signal input
rlabel metal2 s 47030 103200 47086 104000 6 wbs_adr_i[1]
port 520 nsew signal input
rlabel metal2 s 78586 103200 78642 104000 6 wbs_adr_i[20]
port 521 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 wbs_adr_i[21]
port 522 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 wbs_adr_i[22]
port 523 nsew signal input
rlabel metal3 s 103200 32648 104000 32768 6 wbs_adr_i[23]
port 524 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 wbs_adr_i[24]
port 525 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_adr_i[25]
port 526 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[26]
port 527 nsew signal input
rlabel metal2 s 15474 103200 15530 104000 6 wbs_adr_i[27]
port 528 nsew signal input
rlabel metal3 s 103200 72088 104000 72208 6 wbs_adr_i[28]
port 529 nsew signal input
rlabel metal2 s 92754 103200 92810 104000 6 wbs_adr_i[29]
port 530 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[2]
port 531 nsew signal input
rlabel metal2 s 66350 103200 66406 104000 6 wbs_adr_i[30]
port 532 nsew signal input
rlabel metal3 s 103200 53048 104000 53168 6 wbs_adr_i[31]
port 533 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 wbs_adr_i[3]
port 534 nsew signal input
rlabel metal2 s 64418 103200 64474 104000 6 wbs_adr_i[4]
port 535 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 wbs_adr_i[5]
port 536 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[6]
port 537 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[7]
port 538 nsew signal input
rlabel metal3 s 103200 4088 104000 4208 6 wbs_adr_i[8]
port 539 nsew signal input
rlabel metal3 s 103200 34688 104000 34808 6 wbs_adr_i[9]
port 540 nsew signal input
rlabel metal2 s 16762 103200 16818 104000 6 wbs_cyc_i
port 541 nsew signal input
rlabel metal3 s 103200 103368 104000 103488 6 wbs_dat_i[0]
port 542 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 wbs_dat_i[10]
port 543 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 wbs_dat_i[11]
port 544 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wbs_dat_i[12]
port 545 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[13]
port 546 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[14]
port 547 nsew signal input
rlabel metal3 s 103200 62568 104000 62688 6 wbs_dat_i[15]
port 548 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_i[16]
port 549 nsew signal input
rlabel metal2 s 58622 103200 58678 104000 6 wbs_dat_i[17]
port 550 nsew signal input
rlabel metal2 s 85026 103200 85082 104000 6 wbs_dat_i[18]
port 551 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 wbs_dat_i[19]
port 552 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[1]
port 553 nsew signal input
rlabel metal3 s 103200 70048 104000 70168 6 wbs_dat_i[20]
port 554 nsew signal input
rlabel metal2 s 88890 103200 88946 104000 6 wbs_dat_i[21]
port 555 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 wbs_dat_i[22]
port 556 nsew signal input
rlabel metal3 s 103200 89768 104000 89888 6 wbs_dat_i[23]
port 557 nsew signal input
rlabel metal3 s 103200 38088 104000 38208 6 wbs_dat_i[24]
port 558 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wbs_dat_i[25]
port 559 nsew signal input
rlabel metal2 s 77942 103200 77998 104000 6 wbs_dat_i[26]
port 560 nsew signal input
rlabel metal2 s 14830 103200 14886 104000 6 wbs_dat_i[27]
port 561 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[28]
port 562 nsew signal input
rlabel metal3 s 103200 68688 104000 68808 6 wbs_dat_i[29]
port 563 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 wbs_dat_i[2]
port 564 nsew signal input
rlabel metal3 s 103200 34008 104000 34128 6 wbs_dat_i[30]
port 565 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 wbs_dat_i[31]
port 566 nsew signal input
rlabel metal3 s 103200 5448 104000 5568 6 wbs_dat_i[3]
port 567 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[4]
port 568 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_i[5]
port 569 nsew signal input
rlabel metal3 s 103200 48968 104000 49088 6 wbs_dat_i[6]
port 570 nsew signal input
rlabel metal2 s 75366 103200 75422 104000 6 wbs_dat_i[7]
port 571 nsew signal input
rlabel metal3 s 103200 99968 104000 100088 6 wbs_dat_i[8]
port 572 nsew signal input
rlabel metal3 s 103200 6128 104000 6248 6 wbs_dat_i[9]
port 573 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[0]
port 574 nsew signal output
rlabel metal3 s 103200 63248 104000 63368 6 wbs_dat_o[10]
port 575 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_o[11]
port 576 nsew signal output
rlabel metal3 s 103200 101328 104000 101448 6 wbs_dat_o[12]
port 577 nsew signal output
rlabel metal2 s 72146 103200 72202 104000 6 wbs_dat_o[13]
port 578 nsew signal output
rlabel metal3 s 103200 12248 104000 12368 6 wbs_dat_o[14]
port 579 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 wbs_dat_o[15]
port 580 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 wbs_dat_o[16]
port 581 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 wbs_dat_o[17]
port 582 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 wbs_dat_o[18]
port 583 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 584 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 wbs_dat_o[1]
port 585 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 wbs_dat_o[20]
port 586 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 wbs_dat_o[21]
port 587 nsew signal output
rlabel metal2 s 25778 103200 25834 104000 6 wbs_dat_o[22]
port 588 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 wbs_dat_o[23]
port 589 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o[24]
port 590 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_o[25]
port 591 nsew signal output
rlabel metal2 s 51538 103200 51594 104000 6 wbs_dat_o[26]
port 592 nsew signal output
rlabel metal2 s 28354 103200 28410 104000 6 wbs_dat_o[27]
port 593 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_o[28]
port 594 nsew signal output
rlabel metal2 s 69570 103200 69626 104000 6 wbs_dat_o[29]
port 595 nsew signal output
rlabel metal3 s 103200 28568 104000 28688 6 wbs_dat_o[2]
port 596 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 wbs_dat_o[30]
port 597 nsew signal output
rlabel metal3 s 103200 81608 104000 81728 6 wbs_dat_o[31]
port 598 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[3]
port 599 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[4]
port 600 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_o[5]
port 601 nsew signal output
rlabel metal3 s 103200 77528 104000 77648 6 wbs_dat_o[6]
port 602 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_o[7]
port 603 nsew signal output
rlabel metal2 s 67638 103200 67694 104000 6 wbs_dat_o[8]
port 604 nsew signal output
rlabel metal2 s 66994 103200 67050 104000 6 wbs_dat_o[9]
port 605 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 wbs_sel_i[0]
port 606 nsew signal input
rlabel metal2 s 12254 103200 12310 104000 6 wbs_sel_i[1]
port 607 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 wbs_sel_i[2]
port 608 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 wbs_sel_i[3]
port 609 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 wbs_stb_i
port 610 nsew signal input
rlabel metal3 s 103200 49648 104000 49768 6 wbs_we_i
port 611 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 104000 104000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5551686
string GDS_FILE /home/marwan/spm_ip/openlane/spm/runs/2023-03-22-16-52-58/results/signoff/spm.magic.gds
string GDS_START 356156
<< end >>

