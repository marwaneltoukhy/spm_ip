magic
tech sky130A
magscale 1 2
timestamp 1679477535
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 14 892 119218 119332
<< metal2 >>
rect 18 119200 74 120000
rect 662 119200 718 120000
rect 1306 119200 1362 120000
rect 2594 119200 2650 120000
rect 3238 119200 3294 120000
rect 3882 119200 3938 120000
rect 4526 119200 4582 120000
rect 5170 119200 5226 120000
rect 6458 119200 6514 120000
rect 7102 119200 7158 120000
rect 7746 119200 7802 120000
rect 8390 119200 8446 120000
rect 9034 119200 9090 120000
rect 10322 119200 10378 120000
rect 10966 119200 11022 120000
rect 11610 119200 11666 120000
rect 12254 119200 12310 120000
rect 12898 119200 12954 120000
rect 14186 119200 14242 120000
rect 14830 119200 14886 120000
rect 15474 119200 15530 120000
rect 16118 119200 16174 120000
rect 16762 119200 16818 120000
rect 18050 119200 18106 120000
rect 18694 119200 18750 120000
rect 19338 119200 19394 120000
rect 19982 119200 20038 120000
rect 20626 119200 20682 120000
rect 21914 119200 21970 120000
rect 22558 119200 22614 120000
rect 23202 119200 23258 120000
rect 23846 119200 23902 120000
rect 24490 119200 24546 120000
rect 25778 119200 25834 120000
rect 26422 119200 26478 120000
rect 27066 119200 27122 120000
rect 27710 119200 27766 120000
rect 28354 119200 28410 120000
rect 29642 119200 29698 120000
rect 30286 119200 30342 120000
rect 30930 119200 30986 120000
rect 31574 119200 31630 120000
rect 32218 119200 32274 120000
rect 33506 119200 33562 120000
rect 34150 119200 34206 120000
rect 34794 119200 34850 120000
rect 35438 119200 35494 120000
rect 36082 119200 36138 120000
rect 37370 119200 37426 120000
rect 38014 119200 38070 120000
rect 38658 119200 38714 120000
rect 39302 119200 39358 120000
rect 39946 119200 40002 120000
rect 41234 119200 41290 120000
rect 41878 119200 41934 120000
rect 42522 119200 42578 120000
rect 43166 119200 43222 120000
rect 43810 119200 43866 120000
rect 45098 119200 45154 120000
rect 45742 119200 45798 120000
rect 46386 119200 46442 120000
rect 47030 119200 47086 120000
rect 47674 119200 47730 120000
rect 48962 119200 49018 120000
rect 49606 119200 49662 120000
rect 50250 119200 50306 120000
rect 50894 119200 50950 120000
rect 51538 119200 51594 120000
rect 52826 119200 52882 120000
rect 53470 119200 53526 120000
rect 54114 119200 54170 120000
rect 54758 119200 54814 120000
rect 55402 119200 55458 120000
rect 56690 119200 56746 120000
rect 57334 119200 57390 120000
rect 57978 119200 58034 120000
rect 58622 119200 58678 120000
rect 59266 119200 59322 120000
rect 60554 119200 60610 120000
rect 61198 119200 61254 120000
rect 61842 119200 61898 120000
rect 62486 119200 62542 120000
rect 63130 119200 63186 120000
rect 64418 119200 64474 120000
rect 65062 119200 65118 120000
rect 65706 119200 65762 120000
rect 66350 119200 66406 120000
rect 66994 119200 67050 120000
rect 68282 119200 68338 120000
rect 68926 119200 68982 120000
rect 69570 119200 69626 120000
rect 70214 119200 70270 120000
rect 70858 119200 70914 120000
rect 72146 119200 72202 120000
rect 72790 119200 72846 120000
rect 73434 119200 73490 120000
rect 74078 119200 74134 120000
rect 74722 119200 74778 120000
rect 76010 119200 76066 120000
rect 76654 119200 76710 120000
rect 77298 119200 77354 120000
rect 77942 119200 77998 120000
rect 78586 119200 78642 120000
rect 79874 119200 79930 120000
rect 80518 119200 80574 120000
rect 81162 119200 81218 120000
rect 81806 119200 81862 120000
rect 82450 119200 82506 120000
rect 83738 119200 83794 120000
rect 84382 119200 84438 120000
rect 85026 119200 85082 120000
rect 85670 119200 85726 120000
rect 86314 119200 86370 120000
rect 87602 119200 87658 120000
rect 88246 119200 88302 120000
rect 88890 119200 88946 120000
rect 89534 119200 89590 120000
rect 90178 119200 90234 120000
rect 91466 119200 91522 120000
rect 92110 119200 92166 120000
rect 92754 119200 92810 120000
rect 93398 119200 93454 120000
rect 94042 119200 94098 120000
rect 95330 119200 95386 120000
rect 95974 119200 96030 120000
rect 96618 119200 96674 120000
rect 97262 119200 97318 120000
rect 97906 119200 97962 120000
rect 99194 119200 99250 120000
rect 99838 119200 99894 120000
rect 100482 119200 100538 120000
rect 101126 119200 101182 120000
rect 101770 119200 101826 120000
rect 103058 119200 103114 120000
rect 103702 119200 103758 120000
rect 104346 119200 104402 120000
rect 104990 119200 105046 120000
rect 105634 119200 105690 120000
rect 106922 119200 106978 120000
rect 107566 119200 107622 120000
rect 108210 119200 108266 120000
rect 108854 119200 108910 120000
rect 109498 119200 109554 120000
rect 110786 119200 110842 120000
rect 111430 119200 111486 120000
rect 112074 119200 112130 120000
rect 112718 119200 112774 120000
rect 113362 119200 113418 120000
rect 114650 119200 114706 120000
rect 115294 119200 115350 120000
rect 115938 119200 115994 120000
rect 116582 119200 116638 120000
rect 117226 119200 117282 120000
rect 118514 119200 118570 120000
rect 119158 119200 119214 120000
rect 119802 119200 119858 120000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103702 0 103758 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112718 0 112774 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 114650 0 114706 800
rect 115294 0 115350 800
rect 116582 0 116638 800
rect 117226 0 117282 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119158 0 119214 800
<< obsm2 >>
rect 130 119144 606 119785
rect 774 119144 1250 119785
rect 1418 119144 2538 119785
rect 2706 119144 3182 119785
rect 3350 119144 3826 119785
rect 3994 119144 4470 119785
rect 4638 119144 5114 119785
rect 5282 119144 6402 119785
rect 6570 119144 7046 119785
rect 7214 119144 7690 119785
rect 7858 119144 8334 119785
rect 8502 119144 8978 119785
rect 9146 119144 10266 119785
rect 10434 119144 10910 119785
rect 11078 119144 11554 119785
rect 11722 119144 12198 119785
rect 12366 119144 12842 119785
rect 13010 119144 14130 119785
rect 14298 119144 14774 119785
rect 14942 119144 15418 119785
rect 15586 119144 16062 119785
rect 16230 119144 16706 119785
rect 16874 119144 17994 119785
rect 18162 119144 18638 119785
rect 18806 119144 19282 119785
rect 19450 119144 19926 119785
rect 20094 119144 20570 119785
rect 20738 119144 21858 119785
rect 22026 119144 22502 119785
rect 22670 119144 23146 119785
rect 23314 119144 23790 119785
rect 23958 119144 24434 119785
rect 24602 119144 25722 119785
rect 25890 119144 26366 119785
rect 26534 119144 27010 119785
rect 27178 119144 27654 119785
rect 27822 119144 28298 119785
rect 28466 119144 29586 119785
rect 29754 119144 30230 119785
rect 30398 119144 30874 119785
rect 31042 119144 31518 119785
rect 31686 119144 32162 119785
rect 32330 119144 33450 119785
rect 33618 119144 34094 119785
rect 34262 119144 34738 119785
rect 34906 119144 35382 119785
rect 35550 119144 36026 119785
rect 36194 119144 37314 119785
rect 37482 119144 37958 119785
rect 38126 119144 38602 119785
rect 38770 119144 39246 119785
rect 39414 119144 39890 119785
rect 40058 119144 41178 119785
rect 41346 119144 41822 119785
rect 41990 119144 42466 119785
rect 42634 119144 43110 119785
rect 43278 119144 43754 119785
rect 43922 119144 45042 119785
rect 45210 119144 45686 119785
rect 45854 119144 46330 119785
rect 46498 119144 46974 119785
rect 47142 119144 47618 119785
rect 47786 119144 48906 119785
rect 49074 119144 49550 119785
rect 49718 119144 50194 119785
rect 50362 119144 50838 119785
rect 51006 119144 51482 119785
rect 51650 119144 52770 119785
rect 52938 119144 53414 119785
rect 53582 119144 54058 119785
rect 54226 119144 54702 119785
rect 54870 119144 55346 119785
rect 55514 119144 56634 119785
rect 56802 119144 57278 119785
rect 57446 119144 57922 119785
rect 58090 119144 58566 119785
rect 58734 119144 59210 119785
rect 59378 119144 60498 119785
rect 60666 119144 61142 119785
rect 61310 119144 61786 119785
rect 61954 119144 62430 119785
rect 62598 119144 63074 119785
rect 63242 119144 64362 119785
rect 64530 119144 65006 119785
rect 65174 119144 65650 119785
rect 65818 119144 66294 119785
rect 66462 119144 66938 119785
rect 67106 119144 68226 119785
rect 68394 119144 68870 119785
rect 69038 119144 69514 119785
rect 69682 119144 70158 119785
rect 70326 119144 70802 119785
rect 70970 119144 72090 119785
rect 72258 119144 72734 119785
rect 72902 119144 73378 119785
rect 73546 119144 74022 119785
rect 74190 119144 74666 119785
rect 74834 119144 75954 119785
rect 76122 119144 76598 119785
rect 76766 119144 77242 119785
rect 77410 119144 77886 119785
rect 78054 119144 78530 119785
rect 78698 119144 79818 119785
rect 79986 119144 80462 119785
rect 80630 119144 81106 119785
rect 81274 119144 81750 119785
rect 81918 119144 82394 119785
rect 82562 119144 83682 119785
rect 83850 119144 84326 119785
rect 84494 119144 84970 119785
rect 85138 119144 85614 119785
rect 85782 119144 86258 119785
rect 86426 119144 87546 119785
rect 87714 119144 88190 119785
rect 88358 119144 88834 119785
rect 89002 119144 89478 119785
rect 89646 119144 90122 119785
rect 90290 119144 91410 119785
rect 91578 119144 92054 119785
rect 92222 119144 92698 119785
rect 92866 119144 93342 119785
rect 93510 119144 93986 119785
rect 94154 119144 95274 119785
rect 95442 119144 95918 119785
rect 96086 119144 96562 119785
rect 96730 119144 97206 119785
rect 97374 119144 97850 119785
rect 98018 119144 99138 119785
rect 99306 119144 99782 119785
rect 99950 119144 100426 119785
rect 100594 119144 101070 119785
rect 101238 119144 101714 119785
rect 101882 119144 103002 119785
rect 103170 119144 103646 119785
rect 103814 119144 104290 119785
rect 104458 119144 104934 119785
rect 105102 119144 105578 119785
rect 105746 119144 106866 119785
rect 107034 119144 107510 119785
rect 107678 119144 108154 119785
rect 108322 119144 108798 119785
rect 108966 119144 109442 119785
rect 109610 119144 110730 119785
rect 110898 119144 111374 119785
rect 111542 119144 112018 119785
rect 112186 119144 112662 119785
rect 112830 119144 113306 119785
rect 113474 119144 114594 119785
rect 114762 119144 115238 119785
rect 115406 119144 115882 119785
rect 116050 119144 116526 119785
rect 116694 119144 117170 119785
rect 117338 119144 118458 119785
rect 118626 119144 119102 119785
rect 20 856 119212 119144
rect 130 711 606 856
rect 774 711 1250 856
rect 1418 711 1894 856
rect 2062 711 2538 856
rect 2706 711 3182 856
rect 3350 711 4470 856
rect 4638 711 5114 856
rect 5282 711 5758 856
rect 5926 711 6402 856
rect 6570 711 7046 856
rect 7214 711 8334 856
rect 8502 711 8978 856
rect 9146 711 9622 856
rect 9790 711 10266 856
rect 10434 711 10910 856
rect 11078 711 12198 856
rect 12366 711 12842 856
rect 13010 711 13486 856
rect 13654 711 14130 856
rect 14298 711 14774 856
rect 14942 711 16062 856
rect 16230 711 16706 856
rect 16874 711 17350 856
rect 17518 711 17994 856
rect 18162 711 18638 856
rect 18806 711 19926 856
rect 20094 711 20570 856
rect 20738 711 21214 856
rect 21382 711 21858 856
rect 22026 711 22502 856
rect 22670 711 23790 856
rect 23958 711 24434 856
rect 24602 711 25078 856
rect 25246 711 25722 856
rect 25890 711 26366 856
rect 26534 711 27654 856
rect 27822 711 28298 856
rect 28466 711 28942 856
rect 29110 711 29586 856
rect 29754 711 30230 856
rect 30398 711 31518 856
rect 31686 711 32162 856
rect 32330 711 32806 856
rect 32974 711 33450 856
rect 33618 711 34094 856
rect 34262 711 35382 856
rect 35550 711 36026 856
rect 36194 711 36670 856
rect 36838 711 37314 856
rect 37482 711 37958 856
rect 38126 711 39246 856
rect 39414 711 39890 856
rect 40058 711 40534 856
rect 40702 711 41178 856
rect 41346 711 41822 856
rect 41990 711 43110 856
rect 43278 711 43754 856
rect 43922 711 44398 856
rect 44566 711 45042 856
rect 45210 711 45686 856
rect 45854 711 46974 856
rect 47142 711 47618 856
rect 47786 711 48262 856
rect 48430 711 48906 856
rect 49074 711 49550 856
rect 49718 711 50838 856
rect 51006 711 51482 856
rect 51650 711 52126 856
rect 52294 711 52770 856
rect 52938 711 53414 856
rect 53582 711 54702 856
rect 54870 711 55346 856
rect 55514 711 55990 856
rect 56158 711 56634 856
rect 56802 711 57278 856
rect 57446 711 58566 856
rect 58734 711 59210 856
rect 59378 711 59854 856
rect 60022 711 60498 856
rect 60666 711 61142 856
rect 61310 711 62430 856
rect 62598 711 63074 856
rect 63242 711 63718 856
rect 63886 711 64362 856
rect 64530 711 65006 856
rect 65174 711 66294 856
rect 66462 711 66938 856
rect 67106 711 67582 856
rect 67750 711 68226 856
rect 68394 711 68870 856
rect 69038 711 70158 856
rect 70326 711 70802 856
rect 70970 711 71446 856
rect 71614 711 72090 856
rect 72258 711 72734 856
rect 72902 711 74022 856
rect 74190 711 74666 856
rect 74834 711 75310 856
rect 75478 711 75954 856
rect 76122 711 76598 856
rect 76766 711 77886 856
rect 78054 711 78530 856
rect 78698 711 79174 856
rect 79342 711 79818 856
rect 79986 711 80462 856
rect 80630 711 81750 856
rect 81918 711 82394 856
rect 82562 711 83038 856
rect 83206 711 83682 856
rect 83850 711 84326 856
rect 84494 711 85614 856
rect 85782 711 86258 856
rect 86426 711 86902 856
rect 87070 711 87546 856
rect 87714 711 88190 856
rect 88358 711 89478 856
rect 89646 711 90122 856
rect 90290 711 90766 856
rect 90934 711 91410 856
rect 91578 711 92054 856
rect 92222 711 93342 856
rect 93510 711 93986 856
rect 94154 711 94630 856
rect 94798 711 95274 856
rect 95442 711 95918 856
rect 96086 711 97206 856
rect 97374 711 97850 856
rect 98018 711 98494 856
rect 98662 711 99138 856
rect 99306 711 99782 856
rect 99950 711 101070 856
rect 101238 711 101714 856
rect 101882 711 102358 856
rect 102526 711 103002 856
rect 103170 711 103646 856
rect 103814 711 104934 856
rect 105102 711 105578 856
rect 105746 711 106222 856
rect 106390 711 106866 856
rect 107034 711 107510 856
rect 107678 711 108798 856
rect 108966 711 109442 856
rect 109610 711 110086 856
rect 110254 711 110730 856
rect 110898 711 111374 856
rect 111542 711 112662 856
rect 112830 711 113306 856
rect 113474 711 113950 856
rect 114118 711 114594 856
rect 114762 711 115238 856
rect 115406 711 116526 856
rect 116694 711 117170 856
rect 117338 711 117814 856
rect 117982 711 118458 856
rect 118626 711 119102 856
<< metal3 >>
rect 0 119688 800 119808
rect 119200 119688 120000 119808
rect 0 119008 800 119128
rect 119200 119008 120000 119128
rect 119200 118328 120000 118448
rect 0 117648 800 117768
rect 0 116968 800 117088
rect 119200 116968 120000 117088
rect 0 116288 800 116408
rect 119200 116288 120000 116408
rect 0 115608 800 115728
rect 119200 115608 120000 115728
rect 0 114928 800 115048
rect 119200 114928 120000 115048
rect 119200 114248 120000 114368
rect 0 113568 800 113688
rect 0 112888 800 113008
rect 119200 112888 120000 113008
rect 0 112208 800 112328
rect 119200 112208 120000 112328
rect 0 111528 800 111648
rect 119200 111528 120000 111648
rect 0 110848 800 110968
rect 119200 110848 120000 110968
rect 119200 110168 120000 110288
rect 0 109488 800 109608
rect 0 108808 800 108928
rect 119200 108808 120000 108928
rect 0 108128 800 108248
rect 119200 108128 120000 108248
rect 0 107448 800 107568
rect 119200 107448 120000 107568
rect 0 106768 800 106888
rect 119200 106768 120000 106888
rect 119200 106088 120000 106208
rect 0 105408 800 105528
rect 0 104728 800 104848
rect 119200 104728 120000 104848
rect 0 104048 800 104168
rect 119200 104048 120000 104168
rect 0 103368 800 103488
rect 119200 103368 120000 103488
rect 0 102688 800 102808
rect 119200 102688 120000 102808
rect 119200 102008 120000 102128
rect 0 101328 800 101448
rect 0 100648 800 100768
rect 119200 100648 120000 100768
rect 0 99968 800 100088
rect 119200 99968 120000 100088
rect 0 99288 800 99408
rect 119200 99288 120000 99408
rect 0 98608 800 98728
rect 119200 98608 120000 98728
rect 119200 97928 120000 98048
rect 0 97248 800 97368
rect 0 96568 800 96688
rect 119200 96568 120000 96688
rect 0 95888 800 96008
rect 119200 95888 120000 96008
rect 0 95208 800 95328
rect 119200 95208 120000 95328
rect 0 94528 800 94648
rect 119200 94528 120000 94648
rect 119200 93848 120000 93968
rect 0 93168 800 93288
rect 0 92488 800 92608
rect 119200 92488 120000 92608
rect 0 91808 800 91928
rect 119200 91808 120000 91928
rect 0 91128 800 91248
rect 119200 91128 120000 91248
rect 0 90448 800 90568
rect 119200 90448 120000 90568
rect 119200 89768 120000 89888
rect 0 89088 800 89208
rect 0 88408 800 88528
rect 119200 88408 120000 88528
rect 0 87728 800 87848
rect 119200 87728 120000 87848
rect 0 87048 800 87168
rect 119200 87048 120000 87168
rect 0 86368 800 86488
rect 119200 86368 120000 86488
rect 119200 85688 120000 85808
rect 0 85008 800 85128
rect 0 84328 800 84448
rect 119200 84328 120000 84448
rect 0 83648 800 83768
rect 119200 83648 120000 83768
rect 0 82968 800 83088
rect 119200 82968 120000 83088
rect 0 82288 800 82408
rect 119200 82288 120000 82408
rect 119200 81608 120000 81728
rect 0 80928 800 81048
rect 0 80248 800 80368
rect 119200 80248 120000 80368
rect 0 79568 800 79688
rect 119200 79568 120000 79688
rect 0 78888 800 79008
rect 119200 78888 120000 79008
rect 0 78208 800 78328
rect 119200 78208 120000 78328
rect 119200 77528 120000 77648
rect 0 76848 800 76968
rect 0 76168 800 76288
rect 119200 76168 120000 76288
rect 0 75488 800 75608
rect 119200 75488 120000 75608
rect 0 74808 800 74928
rect 119200 74808 120000 74928
rect 0 74128 800 74248
rect 119200 74128 120000 74248
rect 119200 73448 120000 73568
rect 0 72768 800 72888
rect 0 72088 800 72208
rect 119200 72088 120000 72208
rect 0 71408 800 71528
rect 119200 71408 120000 71528
rect 0 70728 800 70848
rect 119200 70728 120000 70848
rect 0 70048 800 70168
rect 119200 70048 120000 70168
rect 119200 69368 120000 69488
rect 0 68688 800 68808
rect 0 68008 800 68128
rect 119200 68008 120000 68128
rect 0 67328 800 67448
rect 119200 67328 120000 67448
rect 0 66648 800 66768
rect 119200 66648 120000 66768
rect 0 65968 800 66088
rect 119200 65968 120000 66088
rect 119200 65288 120000 65408
rect 0 64608 800 64728
rect 0 63928 800 64048
rect 119200 63928 120000 64048
rect 0 63248 800 63368
rect 119200 63248 120000 63368
rect 0 62568 800 62688
rect 119200 62568 120000 62688
rect 0 61888 800 62008
rect 119200 61888 120000 62008
rect 119200 61208 120000 61328
rect 0 60528 800 60648
rect 0 59848 800 59968
rect 119200 59848 120000 59968
rect 0 59168 800 59288
rect 119200 59168 120000 59288
rect 0 58488 800 58608
rect 119200 58488 120000 58608
rect 0 57808 800 57928
rect 119200 57808 120000 57928
rect 119200 57128 120000 57248
rect 0 56448 800 56568
rect 0 55768 800 55888
rect 119200 55768 120000 55888
rect 0 55088 800 55208
rect 119200 55088 120000 55208
rect 0 54408 800 54528
rect 119200 54408 120000 54528
rect 0 53728 800 53848
rect 119200 53728 120000 53848
rect 119200 53048 120000 53168
rect 0 52368 800 52488
rect 0 51688 800 51808
rect 119200 51688 120000 51808
rect 0 51008 800 51128
rect 119200 51008 120000 51128
rect 0 50328 800 50448
rect 119200 50328 120000 50448
rect 0 49648 800 49768
rect 119200 49648 120000 49768
rect 119200 48968 120000 49088
rect 0 48288 800 48408
rect 0 47608 800 47728
rect 119200 47608 120000 47728
rect 0 46928 800 47048
rect 119200 46928 120000 47048
rect 0 46248 800 46368
rect 119200 46248 120000 46368
rect 0 45568 800 45688
rect 119200 45568 120000 45688
rect 119200 44888 120000 45008
rect 0 44208 800 44328
rect 0 43528 800 43648
rect 119200 43528 120000 43648
rect 0 42848 800 42968
rect 119200 42848 120000 42968
rect 0 42168 800 42288
rect 119200 42168 120000 42288
rect 0 41488 800 41608
rect 119200 41488 120000 41608
rect 119200 40808 120000 40928
rect 0 40128 800 40248
rect 0 39448 800 39568
rect 119200 39448 120000 39568
rect 0 38768 800 38888
rect 119200 38768 120000 38888
rect 0 38088 800 38208
rect 119200 38088 120000 38208
rect 0 37408 800 37528
rect 119200 37408 120000 37528
rect 119200 36728 120000 36848
rect 0 36048 800 36168
rect 0 35368 800 35488
rect 119200 35368 120000 35488
rect 0 34688 800 34808
rect 119200 34688 120000 34808
rect 0 34008 800 34128
rect 119200 34008 120000 34128
rect 0 33328 800 33448
rect 119200 33328 120000 33448
rect 119200 32648 120000 32768
rect 0 31968 800 32088
rect 0 31288 800 31408
rect 119200 31288 120000 31408
rect 0 30608 800 30728
rect 119200 30608 120000 30728
rect 0 29928 800 30048
rect 119200 29928 120000 30048
rect 0 29248 800 29368
rect 119200 29248 120000 29368
rect 119200 28568 120000 28688
rect 0 27888 800 28008
rect 0 27208 800 27328
rect 119200 27208 120000 27328
rect 0 26528 800 26648
rect 119200 26528 120000 26648
rect 0 25848 800 25968
rect 119200 25848 120000 25968
rect 0 25168 800 25288
rect 119200 25168 120000 25288
rect 119200 24488 120000 24608
rect 0 23808 800 23928
rect 0 23128 800 23248
rect 119200 23128 120000 23248
rect 0 22448 800 22568
rect 119200 22448 120000 22568
rect 0 21768 800 21888
rect 119200 21768 120000 21888
rect 0 21088 800 21208
rect 119200 21088 120000 21208
rect 119200 20408 120000 20528
rect 0 19728 800 19848
rect 0 19048 800 19168
rect 119200 19048 120000 19168
rect 0 18368 800 18488
rect 119200 18368 120000 18488
rect 0 17688 800 17808
rect 119200 17688 120000 17808
rect 0 17008 800 17128
rect 119200 17008 120000 17128
rect 119200 16328 120000 16448
rect 0 15648 800 15768
rect 0 14968 800 15088
rect 119200 14968 120000 15088
rect 0 14288 800 14408
rect 119200 14288 120000 14408
rect 0 13608 800 13728
rect 119200 13608 120000 13728
rect 0 12928 800 13048
rect 119200 12928 120000 13048
rect 119200 12248 120000 12368
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 119200 10888 120000 11008
rect 0 10208 800 10328
rect 119200 10208 120000 10328
rect 0 9528 800 9648
rect 119200 9528 120000 9648
rect 0 8848 800 8968
rect 119200 8848 120000 8968
rect 119200 8168 120000 8288
rect 0 7488 800 7608
rect 0 6808 800 6928
rect 119200 6808 120000 6928
rect 0 6128 800 6248
rect 119200 6128 120000 6248
rect 0 5448 800 5568
rect 119200 5448 120000 5568
rect 0 4768 800 4888
rect 119200 4768 120000 4888
rect 119200 4088 120000 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
rect 119200 2728 120000 2848
rect 0 2048 800 2168
rect 119200 2048 120000 2168
rect 0 1368 800 1488
rect 119200 1368 120000 1488
rect 0 688 800 808
rect 119200 688 120000 808
rect 119200 8 120000 128
<< obsm3 >>
rect 880 119608 119120 119781
rect 800 119208 119200 119608
rect 880 118928 119120 119208
rect 800 118528 119200 118928
rect 800 118248 119120 118528
rect 800 117848 119200 118248
rect 880 117568 119200 117848
rect 800 117168 119200 117568
rect 880 116888 119120 117168
rect 800 116488 119200 116888
rect 880 116208 119120 116488
rect 800 115808 119200 116208
rect 880 115528 119120 115808
rect 800 115128 119200 115528
rect 880 114848 119120 115128
rect 800 114448 119200 114848
rect 800 114168 119120 114448
rect 800 113768 119200 114168
rect 880 113488 119200 113768
rect 800 113088 119200 113488
rect 880 112808 119120 113088
rect 800 112408 119200 112808
rect 880 112128 119120 112408
rect 800 111728 119200 112128
rect 880 111448 119120 111728
rect 800 111048 119200 111448
rect 880 110768 119120 111048
rect 800 110368 119200 110768
rect 800 110088 119120 110368
rect 800 109688 119200 110088
rect 880 109408 119200 109688
rect 800 109008 119200 109408
rect 880 108728 119120 109008
rect 800 108328 119200 108728
rect 880 108048 119120 108328
rect 800 107648 119200 108048
rect 880 107368 119120 107648
rect 800 106968 119200 107368
rect 880 106688 119120 106968
rect 800 106288 119200 106688
rect 800 106008 119120 106288
rect 800 105608 119200 106008
rect 880 105328 119200 105608
rect 800 104928 119200 105328
rect 880 104648 119120 104928
rect 800 104248 119200 104648
rect 880 103968 119120 104248
rect 800 103568 119200 103968
rect 880 103288 119120 103568
rect 800 102888 119200 103288
rect 880 102608 119120 102888
rect 800 102208 119200 102608
rect 800 101928 119120 102208
rect 800 101528 119200 101928
rect 880 101248 119200 101528
rect 800 100848 119200 101248
rect 880 100568 119120 100848
rect 800 100168 119200 100568
rect 880 99888 119120 100168
rect 800 99488 119200 99888
rect 880 99208 119120 99488
rect 800 98808 119200 99208
rect 880 98528 119120 98808
rect 800 98128 119200 98528
rect 800 97848 119120 98128
rect 800 97448 119200 97848
rect 880 97168 119200 97448
rect 800 96768 119200 97168
rect 880 96488 119120 96768
rect 800 96088 119200 96488
rect 880 95808 119120 96088
rect 800 95408 119200 95808
rect 880 95128 119120 95408
rect 800 94728 119200 95128
rect 880 94448 119120 94728
rect 800 94048 119200 94448
rect 800 93768 119120 94048
rect 800 93368 119200 93768
rect 880 93088 119200 93368
rect 800 92688 119200 93088
rect 880 92408 119120 92688
rect 800 92008 119200 92408
rect 880 91728 119120 92008
rect 800 91328 119200 91728
rect 880 91048 119120 91328
rect 800 90648 119200 91048
rect 880 90368 119120 90648
rect 800 89968 119200 90368
rect 800 89688 119120 89968
rect 800 89288 119200 89688
rect 880 89008 119200 89288
rect 800 88608 119200 89008
rect 880 88328 119120 88608
rect 800 87928 119200 88328
rect 880 87648 119120 87928
rect 800 87248 119200 87648
rect 880 86968 119120 87248
rect 800 86568 119200 86968
rect 880 86288 119120 86568
rect 800 85888 119200 86288
rect 800 85608 119120 85888
rect 800 85208 119200 85608
rect 880 84928 119200 85208
rect 800 84528 119200 84928
rect 880 84248 119120 84528
rect 800 83848 119200 84248
rect 880 83568 119120 83848
rect 800 83168 119200 83568
rect 880 82888 119120 83168
rect 800 82488 119200 82888
rect 880 82208 119120 82488
rect 800 81808 119200 82208
rect 800 81528 119120 81808
rect 800 81128 119200 81528
rect 880 80848 119200 81128
rect 800 80448 119200 80848
rect 880 80168 119120 80448
rect 800 79768 119200 80168
rect 880 79488 119120 79768
rect 800 79088 119200 79488
rect 880 78808 119120 79088
rect 800 78408 119200 78808
rect 880 78128 119120 78408
rect 800 77728 119200 78128
rect 800 77448 119120 77728
rect 800 77048 119200 77448
rect 880 76768 119200 77048
rect 800 76368 119200 76768
rect 880 76088 119120 76368
rect 800 75688 119200 76088
rect 880 75408 119120 75688
rect 800 75008 119200 75408
rect 880 74728 119120 75008
rect 800 74328 119200 74728
rect 880 74048 119120 74328
rect 800 73648 119200 74048
rect 800 73368 119120 73648
rect 800 72968 119200 73368
rect 880 72688 119200 72968
rect 800 72288 119200 72688
rect 880 72008 119120 72288
rect 800 71608 119200 72008
rect 880 71328 119120 71608
rect 800 70928 119200 71328
rect 880 70648 119120 70928
rect 800 70248 119200 70648
rect 880 69968 119120 70248
rect 800 69568 119200 69968
rect 800 69288 119120 69568
rect 800 68888 119200 69288
rect 880 68608 119200 68888
rect 800 68208 119200 68608
rect 880 67928 119120 68208
rect 800 67528 119200 67928
rect 880 67248 119120 67528
rect 800 66848 119200 67248
rect 880 66568 119120 66848
rect 800 66168 119200 66568
rect 880 65888 119120 66168
rect 800 65488 119200 65888
rect 800 65208 119120 65488
rect 800 64808 119200 65208
rect 880 64528 119200 64808
rect 800 64128 119200 64528
rect 880 63848 119120 64128
rect 800 63448 119200 63848
rect 880 63168 119120 63448
rect 800 62768 119200 63168
rect 880 62488 119120 62768
rect 800 62088 119200 62488
rect 880 61808 119120 62088
rect 800 61408 119200 61808
rect 800 61128 119120 61408
rect 800 60728 119200 61128
rect 880 60448 119200 60728
rect 800 60048 119200 60448
rect 880 59768 119120 60048
rect 800 59368 119200 59768
rect 880 59088 119120 59368
rect 800 58688 119200 59088
rect 880 58408 119120 58688
rect 800 58008 119200 58408
rect 880 57728 119120 58008
rect 800 57328 119200 57728
rect 800 57048 119120 57328
rect 800 56648 119200 57048
rect 880 56368 119200 56648
rect 800 55968 119200 56368
rect 880 55688 119120 55968
rect 800 55288 119200 55688
rect 880 55008 119120 55288
rect 800 54608 119200 55008
rect 880 54328 119120 54608
rect 800 53928 119200 54328
rect 880 53648 119120 53928
rect 800 53248 119200 53648
rect 800 52968 119120 53248
rect 800 52568 119200 52968
rect 880 52288 119200 52568
rect 800 51888 119200 52288
rect 880 51608 119120 51888
rect 800 51208 119200 51608
rect 880 50928 119120 51208
rect 800 50528 119200 50928
rect 880 50248 119120 50528
rect 800 49848 119200 50248
rect 880 49568 119120 49848
rect 800 49168 119200 49568
rect 800 48888 119120 49168
rect 800 48488 119200 48888
rect 880 48208 119200 48488
rect 800 47808 119200 48208
rect 880 47528 119120 47808
rect 800 47128 119200 47528
rect 880 46848 119120 47128
rect 800 46448 119200 46848
rect 880 46168 119120 46448
rect 800 45768 119200 46168
rect 880 45488 119120 45768
rect 800 45088 119200 45488
rect 800 44808 119120 45088
rect 800 44408 119200 44808
rect 880 44128 119200 44408
rect 800 43728 119200 44128
rect 880 43448 119120 43728
rect 800 43048 119200 43448
rect 880 42768 119120 43048
rect 800 42368 119200 42768
rect 880 42088 119120 42368
rect 800 41688 119200 42088
rect 880 41408 119120 41688
rect 800 41008 119200 41408
rect 800 40728 119120 41008
rect 800 40328 119200 40728
rect 880 40048 119200 40328
rect 800 39648 119200 40048
rect 880 39368 119120 39648
rect 800 38968 119200 39368
rect 880 38688 119120 38968
rect 800 38288 119200 38688
rect 880 38008 119120 38288
rect 800 37608 119200 38008
rect 880 37328 119120 37608
rect 800 36928 119200 37328
rect 800 36648 119120 36928
rect 800 36248 119200 36648
rect 880 35968 119200 36248
rect 800 35568 119200 35968
rect 880 35288 119120 35568
rect 800 34888 119200 35288
rect 880 34608 119120 34888
rect 800 34208 119200 34608
rect 880 33928 119120 34208
rect 800 33528 119200 33928
rect 880 33248 119120 33528
rect 800 32848 119200 33248
rect 800 32568 119120 32848
rect 800 32168 119200 32568
rect 880 31888 119200 32168
rect 800 31488 119200 31888
rect 880 31208 119120 31488
rect 800 30808 119200 31208
rect 880 30528 119120 30808
rect 800 30128 119200 30528
rect 880 29848 119120 30128
rect 800 29448 119200 29848
rect 880 29168 119120 29448
rect 800 28768 119200 29168
rect 800 28488 119120 28768
rect 800 28088 119200 28488
rect 880 27808 119200 28088
rect 800 27408 119200 27808
rect 880 27128 119120 27408
rect 800 26728 119200 27128
rect 880 26448 119120 26728
rect 800 26048 119200 26448
rect 880 25768 119120 26048
rect 800 25368 119200 25768
rect 880 25088 119120 25368
rect 800 24688 119200 25088
rect 800 24408 119120 24688
rect 800 24008 119200 24408
rect 880 23728 119200 24008
rect 800 23328 119200 23728
rect 880 23048 119120 23328
rect 800 22648 119200 23048
rect 880 22368 119120 22648
rect 800 21968 119200 22368
rect 880 21688 119120 21968
rect 800 21288 119200 21688
rect 880 21008 119120 21288
rect 800 20608 119200 21008
rect 800 20328 119120 20608
rect 800 19928 119200 20328
rect 880 19648 119200 19928
rect 800 19248 119200 19648
rect 880 18968 119120 19248
rect 800 18568 119200 18968
rect 880 18288 119120 18568
rect 800 17888 119200 18288
rect 880 17608 119120 17888
rect 800 17208 119200 17608
rect 880 16928 119120 17208
rect 800 16528 119200 16928
rect 800 16248 119120 16528
rect 800 15848 119200 16248
rect 880 15568 119200 15848
rect 800 15168 119200 15568
rect 880 14888 119120 15168
rect 800 14488 119200 14888
rect 880 14208 119120 14488
rect 800 13808 119200 14208
rect 880 13528 119120 13808
rect 800 13128 119200 13528
rect 880 12848 119120 13128
rect 800 12448 119200 12848
rect 800 12168 119120 12448
rect 800 11768 119200 12168
rect 880 11488 119200 11768
rect 800 11088 119200 11488
rect 880 10808 119120 11088
rect 800 10408 119200 10808
rect 880 10128 119120 10408
rect 800 9728 119200 10128
rect 880 9448 119120 9728
rect 800 9048 119200 9448
rect 880 8768 119120 9048
rect 800 8368 119200 8768
rect 800 8088 119120 8368
rect 800 7688 119200 8088
rect 880 7408 119200 7688
rect 800 7008 119200 7408
rect 880 6728 119120 7008
rect 800 6328 119200 6728
rect 880 6048 119120 6328
rect 800 5648 119200 6048
rect 880 5368 119120 5648
rect 800 4968 119200 5368
rect 880 4688 119120 4968
rect 800 4288 119200 4688
rect 800 4008 119120 4288
rect 800 3608 119200 4008
rect 880 3328 119200 3608
rect 800 2928 119200 3328
rect 880 2648 119120 2928
rect 800 2248 119200 2648
rect 880 1968 119120 2248
rect 800 1568 119200 1968
rect 880 1288 119120 1568
rect 800 888 119200 1288
rect 880 715 119120 888
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2128 5188 117552
rect 5528 2128 5848 117552
rect 6188 2128 6508 117552
rect 34928 2128 35248 117552
rect 35588 2128 35908 117552
rect 36248 2128 36568 117552
rect 36908 2128 37228 117552
rect 65648 2128 65968 117552
rect 66308 2128 66628 117552
rect 66968 2128 67288 117552
rect 67628 2128 67948 117552
rect 96368 2128 96688 117552
rect 97028 2128 97348 117552
rect 97688 2128 98008 117552
rect 98348 2128 98668 117552
<< obsm4 >>
rect 77155 2347 82557 61029
<< metal5 >>
rect 1056 99234 118912 99554
rect 1056 98574 118912 98894
rect 1056 97914 118912 98234
rect 1056 97254 118912 97574
rect 1056 68598 118912 68918
rect 1056 67938 118912 68258
rect 1056 67278 118912 67598
rect 1056 66618 118912 66938
rect 1056 37962 118912 38282
rect 1056 37302 118912 37622
rect 1056 36642 118912 36962
rect 1056 35982 118912 36302
rect 1056 7326 118912 7646
rect 1056 6666 118912 6986
rect 1056 6006 118912 6326
rect 1056 5346 118912 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 118912 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 118912 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 118912 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 97914 118912 98234 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 118912 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 118912 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 118912 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 118912 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 114650 0 114706 800 6 io_in[0]
port 3 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 119200 51688 120000 51808 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 io_in[12]
port 6 nsew signal input
rlabel metal2 s 41234 119200 41290 120000 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 119200 78208 120000 78328 6 io_in[14]
port 8 nsew signal input
rlabel metal2 s 34794 119200 34850 120000 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 119200 114928 120000 115048 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 io_in[18]
port 12 nsew signal input
rlabel metal2 s 45098 119200 45154 120000 6 io_in[19]
port 13 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 io_in[1]
port 14 nsew signal input
rlabel metal2 s 30930 119200 30986 120000 6 io_in[20]
port 15 nsew signal input
rlabel metal2 s 37370 119200 37426 120000 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 119200 88408 120000 88528 6 io_in[24]
port 19 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[25]
port 20 nsew signal input
rlabel metal2 s 76010 119200 76066 120000 6 io_in[26]
port 21 nsew signal input
rlabel metal2 s 33506 119200 33562 120000 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 io_in[28]
port 23 nsew signal input
rlabel metal2 s 54758 119200 54814 120000 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 io_in[2]
port 25 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_in[31]
port 27 nsew signal input
rlabel metal2 s 81806 119200 81862 120000 6 io_in[32]
port 28 nsew signal input
rlabel metal2 s 70214 119200 70270 120000 6 io_in[33]
port 29 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 io_in[34]
port 30 nsew signal input
rlabel metal3 s 119200 78888 120000 79008 6 io_in[35]
port 31 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 io_in[36]
port 32 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 io_in[37]
port 33 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 io_in[3]
port 34 nsew signal input
rlabel metal2 s 113362 119200 113418 120000 6 io_in[4]
port 35 nsew signal input
rlabel metal3 s 119200 12928 120000 13048 6 io_in[5]
port 36 nsew signal input
rlabel metal3 s 119200 70048 120000 70168 6 io_in[6]
port 37 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 io_in[7]
port 38 nsew signal input
rlabel metal2 s 57978 119200 58034 120000 6 io_in[8]
port 39 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 io_in[9]
port 40 nsew signal input
rlabel metal3 s 119200 41488 120000 41608 6 io_oeb[0]
port 41 nsew signal output
rlabel metal3 s 119200 38768 120000 38888 6 io_oeb[10]
port 42 nsew signal output
rlabel metal2 s 72146 119200 72202 120000 6 io_oeb[11]
port 43 nsew signal output
rlabel metal2 s 42522 119200 42578 120000 6 io_oeb[12]
port 44 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 io_oeb[13]
port 45 nsew signal output
rlabel metal2 s 21914 119200 21970 120000 6 io_oeb[14]
port 46 nsew signal output
rlabel metal3 s 119200 42168 120000 42288 6 io_oeb[15]
port 47 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 io_oeb[16]
port 48 nsew signal output
rlabel metal2 s 1306 119200 1362 120000 6 io_oeb[17]
port 49 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 io_oeb[18]
port 50 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 io_oeb[19]
port 51 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 io_oeb[1]
port 52 nsew signal output
rlabel metal2 s 22558 119200 22614 120000 6 io_oeb[20]
port 53 nsew signal output
rlabel metal2 s 82450 119200 82506 120000 6 io_oeb[21]
port 54 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_oeb[22]
port 55 nsew signal output
rlabel metal3 s 119200 47608 120000 47728 6 io_oeb[23]
port 56 nsew signal output
rlabel metal3 s 119200 119008 120000 119128 6 io_oeb[24]
port 57 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 io_oeb[25]
port 58 nsew signal output
rlabel metal2 s 14830 119200 14886 120000 6 io_oeb[26]
port 59 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_oeb[27]
port 60 nsew signal output
rlabel metal2 s 73434 119200 73490 120000 6 io_oeb[28]
port 61 nsew signal output
rlabel metal3 s 119200 87728 120000 87848 6 io_oeb[29]
port 62 nsew signal output
rlabel metal3 s 119200 103368 120000 103488 6 io_oeb[2]
port 63 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 io_oeb[30]
port 64 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 io_oeb[31]
port 65 nsew signal output
rlabel metal2 s 16118 119200 16174 120000 6 io_oeb[32]
port 66 nsew signal output
rlabel metal2 s 6458 119200 6514 120000 6 io_oeb[33]
port 67 nsew signal output
rlabel metal2 s 23202 119200 23258 120000 6 io_oeb[34]
port 68 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 io_oeb[35]
port 69 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 io_oeb[36]
port 70 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 io_oeb[37]
port 71 nsew signal output
rlabel metal2 s 92110 119200 92166 120000 6 io_oeb[3]
port 72 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 io_oeb[4]
port 73 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 io_oeb[5]
port 74 nsew signal output
rlabel metal2 s 86314 119200 86370 120000 6 io_oeb[6]
port 75 nsew signal output
rlabel metal2 s 115938 119200 115994 120000 6 io_oeb[7]
port 76 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 io_oeb[8]
port 77 nsew signal output
rlabel metal2 s 12898 119200 12954 120000 6 io_oeb[9]
port 78 nsew signal output
rlabel metal2 s 18 119200 74 120000 6 io_out[0]
port 79 nsew signal output
rlabel metal2 s 112718 119200 112774 120000 6 io_out[10]
port 80 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 io_out[11]
port 81 nsew signal output
rlabel metal3 s 119200 111528 120000 111648 6 io_out[12]
port 82 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_out[13]
port 83 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 io_out[14]
port 84 nsew signal output
rlabel metal3 s 119200 92488 120000 92608 6 io_out[15]
port 85 nsew signal output
rlabel metal3 s 119200 25848 120000 25968 6 io_out[16]
port 86 nsew signal output
rlabel metal3 s 119200 77528 120000 77648 6 io_out[17]
port 87 nsew signal output
rlabel metal3 s 119200 107448 120000 107568 6 io_out[18]
port 88 nsew signal output
rlabel metal3 s 119200 93848 120000 93968 6 io_out[19]
port 89 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 io_out[1]
port 90 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 io_out[20]
port 91 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 io_out[21]
port 92 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 io_out[22]
port 93 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 io_out[23]
port 94 nsew signal output
rlabel metal3 s 119200 10888 120000 11008 6 io_out[24]
port 95 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 io_out[25]
port 96 nsew signal output
rlabel metal2 s 24490 119200 24546 120000 6 io_out[26]
port 97 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 io_out[27]
port 98 nsew signal output
rlabel metal3 s 119200 65968 120000 66088 6 io_out[28]
port 99 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 io_out[29]
port 100 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 io_out[2]
port 101 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 io_out[30]
port 102 nsew signal output
rlabel metal3 s 119200 106088 120000 106208 6 io_out[31]
port 103 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 io_out[32]
port 104 nsew signal output
rlabel metal3 s 119200 90448 120000 90568 6 io_out[33]
port 105 nsew signal output
rlabel metal2 s 119158 119200 119214 120000 6 io_out[34]
port 106 nsew signal output
rlabel metal3 s 119200 80248 120000 80368 6 io_out[35]
port 107 nsew signal output
rlabel metal2 s 23846 119200 23902 120000 6 io_out[36]
port 108 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 io_out[37]
port 109 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 io_out[3]
port 110 nsew signal output
rlabel metal3 s 119200 9528 120000 9648 6 io_out[4]
port 111 nsew signal output
rlabel metal3 s 119200 74128 120000 74248 6 io_out[5]
port 112 nsew signal output
rlabel metal2 s 61198 119200 61254 120000 6 io_out[6]
port 113 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_out[7]
port 114 nsew signal output
rlabel metal2 s 49606 119200 49662 120000 6 io_out[8]
port 115 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 io_out[9]
port 116 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 irq[0]
port 117 nsew signal output
rlabel metal3 s 119200 46928 120000 47048 6 irq[1]
port 118 nsew signal output
rlabel metal2 s 95330 119200 95386 120000 6 irq[2]
port 119 nsew signal output
rlabel metal3 s 119200 59848 120000 59968 6 la_data_in[0]
port 120 nsew signal input
rlabel metal3 s 119200 32648 120000 32768 6 la_data_in[100]
port 121 nsew signal input
rlabel metal2 s 53470 119200 53526 120000 6 la_data_in[101]
port 122 nsew signal input
rlabel metal2 s 19982 119200 20038 120000 6 la_data_in[102]
port 123 nsew signal input
rlabel metal3 s 119200 110168 120000 110288 6 la_data_in[103]
port 124 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 la_data_in[104]
port 125 nsew signal input
rlabel metal3 s 119200 74808 120000 74928 6 la_data_in[105]
port 126 nsew signal input
rlabel metal3 s 119200 10208 120000 10328 6 la_data_in[106]
port 127 nsew signal input
rlabel metal2 s 65706 119200 65762 120000 6 la_data_in[107]
port 128 nsew signal input
rlabel metal3 s 119200 29928 120000 30048 6 la_data_in[108]
port 129 nsew signal input
rlabel metal2 s 85670 119200 85726 120000 6 la_data_in[109]
port 130 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 la_data_in[10]
port 131 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[110]
port 132 nsew signal input
rlabel metal3 s 119200 75488 120000 75608 6 la_data_in[111]
port 133 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 la_data_in[112]
port 134 nsew signal input
rlabel metal3 s 119200 17008 120000 17128 6 la_data_in[113]
port 135 nsew signal input
rlabel metal2 s 88890 119200 88946 120000 6 la_data_in[114]
port 136 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[115]
port 137 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[116]
port 138 nsew signal input
rlabel metal2 s 48962 119200 49018 120000 6 la_data_in[117]
port 139 nsew signal input
rlabel metal2 s 96618 119200 96674 120000 6 la_data_in[118]
port 140 nsew signal input
rlabel metal3 s 119200 71408 120000 71528 6 la_data_in[119]
port 141 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 la_data_in[11]
port 142 nsew signal input
rlabel metal2 s 81162 119200 81218 120000 6 la_data_in[120]
port 143 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[121]
port 144 nsew signal input
rlabel metal2 s 7102 119200 7158 120000 6 la_data_in[122]
port 145 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[123]
port 146 nsew signal input
rlabel metal2 s 11610 119200 11666 120000 6 la_data_in[124]
port 147 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 la_data_in[125]
port 148 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[126]
port 149 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 la_data_in[127]
port 150 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 la_data_in[12]
port 151 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[13]
port 152 nsew signal input
rlabel metal3 s 119200 86368 120000 86488 6 la_data_in[14]
port 153 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 la_data_in[15]
port 154 nsew signal input
rlabel metal3 s 119200 49648 120000 49768 6 la_data_in[16]
port 155 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 la_data_in[17]
port 156 nsew signal input
rlabel metal3 s 119200 100648 120000 100768 6 la_data_in[18]
port 157 nsew signal input
rlabel metal2 s 91466 119200 91522 120000 6 la_data_in[19]
port 158 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[1]
port 159 nsew signal input
rlabel metal2 s 3238 119200 3294 120000 6 la_data_in[20]
port 160 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_data_in[21]
port 161 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[22]
port 162 nsew signal input
rlabel metal3 s 119200 62568 120000 62688 6 la_data_in[23]
port 163 nsew signal input
rlabel metal3 s 119200 21768 120000 21888 6 la_data_in[24]
port 164 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 la_data_in[25]
port 165 nsew signal input
rlabel metal3 s 119200 95888 120000 96008 6 la_data_in[26]
port 166 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[27]
port 167 nsew signal input
rlabel metal3 s 119200 70728 120000 70848 6 la_data_in[28]
port 168 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[29]
port 169 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[2]
port 170 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[30]
port 171 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 la_data_in[31]
port 172 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[32]
port 173 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[33]
port 174 nsew signal input
rlabel metal2 s 55402 119200 55458 120000 6 la_data_in[34]
port 175 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 la_data_in[35]
port 176 nsew signal input
rlabel metal2 s 94042 119200 94098 120000 6 la_data_in[36]
port 177 nsew signal input
rlabel metal2 s 116582 119200 116638 120000 6 la_data_in[37]
port 178 nsew signal input
rlabel metal3 s 119200 51008 120000 51128 6 la_data_in[38]
port 179 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 la_data_in[39]
port 180 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_data_in[3]
port 181 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_data_in[40]
port 182 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[41]
port 183 nsew signal input
rlabel metal3 s 119200 53728 120000 53848 6 la_data_in[42]
port 184 nsew signal input
rlabel metal3 s 119200 91808 120000 91928 6 la_data_in[43]
port 185 nsew signal input
rlabel metal2 s 39946 119200 40002 120000 6 la_data_in[44]
port 186 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 la_data_in[45]
port 187 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 la_data_in[46]
port 188 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[47]
port 189 nsew signal input
rlabel metal2 s 85026 119200 85082 120000 6 la_data_in[48]
port 190 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[49]
port 191 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[4]
port 192 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 la_data_in[50]
port 193 nsew signal input
rlabel metal2 s 2594 119200 2650 120000 6 la_data_in[51]
port 194 nsew signal input
rlabel metal2 s 114650 119200 114706 120000 6 la_data_in[52]
port 195 nsew signal input
rlabel metal3 s 119200 21088 120000 21208 6 la_data_in[53]
port 196 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 la_data_in[54]
port 197 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[55]
port 198 nsew signal input
rlabel metal2 s 662 0 718 800 6 la_data_in[56]
port 199 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[57]
port 200 nsew signal input
rlabel metal2 s 99838 119200 99894 120000 6 la_data_in[58]
port 201 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[59]
port 202 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 la_data_in[5]
port 203 nsew signal input
rlabel metal2 s 10322 119200 10378 120000 6 la_data_in[60]
port 204 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_data_in[61]
port 205 nsew signal input
rlabel metal3 s 119200 27208 120000 27328 6 la_data_in[62]
port 206 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 la_data_in[63]
port 207 nsew signal input
rlabel metal3 s 119200 112888 120000 113008 6 la_data_in[64]
port 208 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[65]
port 209 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 la_data_in[66]
port 210 nsew signal input
rlabel metal2 s 50250 119200 50306 120000 6 la_data_in[67]
port 211 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la_data_in[68]
port 212 nsew signal input
rlabel metal3 s 119200 87048 120000 87168 6 la_data_in[69]
port 213 nsew signal input
rlabel metal3 s 119200 46248 120000 46368 6 la_data_in[6]
port 214 nsew signal input
rlabel metal3 s 119200 28568 120000 28688 6 la_data_in[70]
port 215 nsew signal input
rlabel metal3 s 119200 20408 120000 20528 6 la_data_in[71]
port 216 nsew signal input
rlabel metal2 s 30286 119200 30342 120000 6 la_data_in[72]
port 217 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_data_in[73]
port 218 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[74]
port 219 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[75]
port 220 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[76]
port 221 nsew signal input
rlabel metal3 s 119200 76168 120000 76288 6 la_data_in[77]
port 222 nsew signal input
rlabel metal3 s 119200 95208 120000 95328 6 la_data_in[78]
port 223 nsew signal input
rlabel metal3 s 119200 31288 120000 31408 6 la_data_in[79]
port 224 nsew signal input
rlabel metal3 s 119200 35368 120000 35488 6 la_data_in[7]
port 225 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[80]
port 226 nsew signal input
rlabel metal3 s 119200 36728 120000 36848 6 la_data_in[81]
port 227 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_data_in[82]
port 228 nsew signal input
rlabel metal2 s 100482 119200 100538 120000 6 la_data_in[83]
port 229 nsew signal input
rlabel metal3 s 0 688 800 808 6 la_data_in[84]
port 230 nsew signal input
rlabel metal2 s 47674 119200 47730 120000 6 la_data_in[85]
port 231 nsew signal input
rlabel metal3 s 119200 84328 120000 84448 6 la_data_in[86]
port 232 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 la_data_in[87]
port 233 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 la_data_in[88]
port 234 nsew signal input
rlabel metal2 s 41878 119200 41934 120000 6 la_data_in[89]
port 235 nsew signal input
rlabel metal2 s 28354 119200 28410 120000 6 la_data_in[8]
port 236 nsew signal input
rlabel metal2 s 69570 119200 69626 120000 6 la_data_in[90]
port 237 nsew signal input
rlabel metal2 s 4526 119200 4582 120000 6 la_data_in[91]
port 238 nsew signal input
rlabel metal3 s 119200 8 120000 128 6 la_data_in[92]
port 239 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[93]
port 240 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[94]
port 241 nsew signal input
rlabel metal3 s 119200 8168 120000 8288 6 la_data_in[95]
port 242 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 la_data_in[96]
port 243 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 la_data_in[97]
port 244 nsew signal input
rlabel metal3 s 119200 55088 120000 55208 6 la_data_in[98]
port 245 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 la_data_in[99]
port 246 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_data_in[9]
port 247 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 la_data_out[0]
port 248 nsew signal output
rlabel metal2 s 111430 119200 111486 120000 6 la_data_out[100]
port 249 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 la_data_out[101]
port 250 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 la_data_out[102]
port 251 nsew signal output
rlabel metal3 s 119200 42848 120000 42968 6 la_data_out[103]
port 252 nsew signal output
rlabel metal3 s 119200 63928 120000 64048 6 la_data_out[104]
port 253 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 la_data_out[105]
port 254 nsew signal output
rlabel metal2 s 27710 119200 27766 120000 6 la_data_out[106]
port 255 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[107]
port 256 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 la_data_out[108]
port 257 nsew signal output
rlabel metal2 s 62486 119200 62542 120000 6 la_data_out[109]
port 258 nsew signal output
rlabel metal2 s 72790 119200 72846 120000 6 la_data_out[10]
port 259 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 la_data_out[110]
port 260 nsew signal output
rlabel metal2 s 88246 119200 88302 120000 6 la_data_out[111]
port 261 nsew signal output
rlabel metal2 s 108854 119200 108910 120000 6 la_data_out[112]
port 262 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 la_data_out[113]
port 263 nsew signal output
rlabel metal2 s 50894 119200 50950 120000 6 la_data_out[114]
port 264 nsew signal output
rlabel metal3 s 119200 104728 120000 104848 6 la_data_out[115]
port 265 nsew signal output
rlabel metal3 s 119200 25168 120000 25288 6 la_data_out[116]
port 266 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 la_data_out[117]
port 267 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[118]
port 268 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 la_data_out[119]
port 269 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[11]
port 270 nsew signal output
rlabel metal3 s 119200 1368 120000 1488 6 la_data_out[120]
port 271 nsew signal output
rlabel metal2 s 20626 119200 20682 120000 6 la_data_out[121]
port 272 nsew signal output
rlabel metal2 s 110786 119200 110842 120000 6 la_data_out[122]
port 273 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 la_data_out[123]
port 274 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la_data_out[124]
port 275 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 la_data_out[125]
port 276 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[126]
port 277 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 la_data_out[127]
port 278 nsew signal output
rlabel metal3 s 119200 106768 120000 106888 6 la_data_out[12]
port 279 nsew signal output
rlabel metal3 s 119200 53048 120000 53168 6 la_data_out[13]
port 280 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 la_data_out[14]
port 281 nsew signal output
rlabel metal3 s 119200 58488 120000 58608 6 la_data_out[15]
port 282 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[16]
port 283 nsew signal output
rlabel metal2 s 10966 119200 11022 120000 6 la_data_out[17]
port 284 nsew signal output
rlabel metal3 s 119200 18368 120000 18488 6 la_data_out[18]
port 285 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 la_data_out[19]
port 286 nsew signal output
rlabel metal2 s 9034 119200 9090 120000 6 la_data_out[1]
port 287 nsew signal output
rlabel metal3 s 119200 116288 120000 116408 6 la_data_out[20]
port 288 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 la_data_out[21]
port 289 nsew signal output
rlabel metal2 s 78586 119200 78642 120000 6 la_data_out[22]
port 290 nsew signal output
rlabel metal3 s 119200 43528 120000 43648 6 la_data_out[23]
port 291 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[24]
port 292 nsew signal output
rlabel metal2 s 66994 119200 67050 120000 6 la_data_out[25]
port 293 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 la_data_out[26]
port 294 nsew signal output
rlabel metal3 s 119200 54408 120000 54528 6 la_data_out[27]
port 295 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out[28]
port 296 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 la_data_out[29]
port 297 nsew signal output
rlabel metal3 s 119200 14968 120000 15088 6 la_data_out[2]
port 298 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[30]
port 299 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 la_data_out[31]
port 300 nsew signal output
rlabel metal2 s 26422 119200 26478 120000 6 la_data_out[32]
port 301 nsew signal output
rlabel metal2 s 68926 119200 68982 120000 6 la_data_out[33]
port 302 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[34]
port 303 nsew signal output
rlabel metal2 s 105634 119200 105690 120000 6 la_data_out[35]
port 304 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 la_data_out[36]
port 305 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 la_data_out[37]
port 306 nsew signal output
rlabel metal2 s 95974 119200 96030 120000 6 la_data_out[38]
port 307 nsew signal output
rlabel metal3 s 119200 30608 120000 30728 6 la_data_out[39]
port 308 nsew signal output
rlabel metal2 s 46386 119200 46442 120000 6 la_data_out[3]
port 309 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 la_data_out[40]
port 310 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[41]
port 311 nsew signal output
rlabel metal2 s 38014 119200 38070 120000 6 la_data_out[42]
port 312 nsew signal output
rlabel metal2 s 34150 119200 34206 120000 6 la_data_out[43]
port 313 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[44]
port 314 nsew signal output
rlabel metal3 s 119200 688 120000 808 6 la_data_out[45]
port 315 nsew signal output
rlabel metal2 s 118514 119200 118570 120000 6 la_data_out[46]
port 316 nsew signal output
rlabel metal2 s 43166 119200 43222 120000 6 la_data_out[47]
port 317 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 la_data_out[48]
port 318 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 la_data_out[49]
port 319 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 la_data_out[4]
port 320 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 la_data_out[50]
port 321 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 la_data_out[51]
port 322 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 la_data_out[52]
port 323 nsew signal output
rlabel metal3 s 119200 59168 120000 59288 6 la_data_out[53]
port 324 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 la_data_out[54]
port 325 nsew signal output
rlabel metal3 s 119200 55768 120000 55888 6 la_data_out[55]
port 326 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 la_data_out[56]
port 327 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[57]
port 328 nsew signal output
rlabel metal2 s 112074 119200 112130 120000 6 la_data_out[58]
port 329 nsew signal output
rlabel metal2 s 92754 119200 92810 120000 6 la_data_out[59]
port 330 nsew signal output
rlabel metal2 s 58622 119200 58678 120000 6 la_data_out[5]
port 331 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 la_data_out[60]
port 332 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[61]
port 333 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 la_data_out[62]
port 334 nsew signal output
rlabel metal3 s 119200 63248 120000 63368 6 la_data_out[63]
port 335 nsew signal output
rlabel metal3 s 119200 24488 120000 24608 6 la_data_out[64]
port 336 nsew signal output
rlabel metal3 s 119200 13608 120000 13728 6 la_data_out[65]
port 337 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[66]
port 338 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[67]
port 339 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[68]
port 340 nsew signal output
rlabel metal2 s 108210 119200 108266 120000 6 la_data_out[69]
port 341 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[6]
port 342 nsew signal output
rlabel metal2 s 47030 119200 47086 120000 6 la_data_out[70]
port 343 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 la_data_out[71]
port 344 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[72]
port 345 nsew signal output
rlabel metal2 s 60554 119200 60610 120000 6 la_data_out[73]
port 346 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[74]
port 347 nsew signal output
rlabel metal3 s 119200 8848 120000 8968 6 la_data_out[75]
port 348 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[76]
port 349 nsew signal output
rlabel metal3 s 119200 23128 120000 23248 6 la_data_out[77]
port 350 nsew signal output
rlabel metal3 s 119200 17688 120000 17808 6 la_data_out[78]
port 351 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[79]
port 352 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 la_data_out[7]
port 353 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 la_data_out[80]
port 354 nsew signal output
rlabel metal2 s 27066 119200 27122 120000 6 la_data_out[81]
port 355 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 la_data_out[82]
port 356 nsew signal output
rlabel metal2 s 18694 119200 18750 120000 6 la_data_out[83]
port 357 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 la_data_out[84]
port 358 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[85]
port 359 nsew signal output
rlabel metal3 s 119200 61208 120000 61328 6 la_data_out[86]
port 360 nsew signal output
rlabel metal2 s 66350 119200 66406 120000 6 la_data_out[87]
port 361 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[88]
port 362 nsew signal output
rlabel metal2 s 63130 119200 63186 120000 6 la_data_out[89]
port 363 nsew signal output
rlabel metal2 s 64418 119200 64474 120000 6 la_data_out[8]
port 364 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[90]
port 365 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[91]
port 366 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 la_data_out[92]
port 367 nsew signal output
rlabel metal2 s 39302 119200 39358 120000 6 la_data_out[93]
port 368 nsew signal output
rlabel metal2 s 51538 119200 51594 120000 6 la_data_out[94]
port 369 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[95]
port 370 nsew signal output
rlabel metal2 s 12254 119200 12310 120000 6 la_data_out[96]
port 371 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 la_data_out[97]
port 372 nsew signal output
rlabel metal2 s 99194 119200 99250 120000 6 la_data_out[98]
port 373 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[99]
port 374 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[9]
port 375 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_oenb[0]
port 376 nsew signal input
rlabel metal3 s 119200 118328 120000 118448 6 la_oenb[100]
port 377 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 la_oenb[101]
port 378 nsew signal input
rlabel metal2 s 101126 119200 101182 120000 6 la_oenb[102]
port 379 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_oenb[103]
port 380 nsew signal input
rlabel metal3 s 119200 68008 120000 68128 6 la_oenb[104]
port 381 nsew signal input
rlabel metal2 s 56690 119200 56746 120000 6 la_oenb[105]
port 382 nsew signal input
rlabel metal2 s 117226 119200 117282 120000 6 la_oenb[106]
port 383 nsew signal input
rlabel metal3 s 119200 66648 120000 66768 6 la_oenb[107]
port 384 nsew signal input
rlabel metal2 s 79874 119200 79930 120000 6 la_oenb[108]
port 385 nsew signal input
rlabel metal2 s 93398 119200 93454 120000 6 la_oenb[109]
port 386 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[10]
port 387 nsew signal input
rlabel metal3 s 119200 91128 120000 91248 6 la_oenb[110]
port 388 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[111]
port 389 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la_oenb[112]
port 390 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la_oenb[113]
port 391 nsew signal input
rlabel metal2 s 70858 119200 70914 120000 6 la_oenb[114]
port 392 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[115]
port 393 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[116]
port 394 nsew signal input
rlabel metal3 s 119200 114248 120000 114368 6 la_oenb[117]
port 395 nsew signal input
rlabel metal3 s 119200 45568 120000 45688 6 la_oenb[118]
port 396 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_oenb[119]
port 397 nsew signal input
rlabel metal3 s 119200 67328 120000 67448 6 la_oenb[11]
port 398 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[120]
port 399 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[121]
port 400 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 la_oenb[122]
port 401 nsew signal input
rlabel metal3 s 119200 99288 120000 99408 6 la_oenb[123]
port 402 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_oenb[124]
port 403 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_oenb[125]
port 404 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[126]
port 405 nsew signal input
rlabel metal3 s 119200 29248 120000 29368 6 la_oenb[127]
port 406 nsew signal input
rlabel metal3 s 119200 82288 120000 82408 6 la_oenb[12]
port 407 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la_oenb[13]
port 408 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_oenb[14]
port 409 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[15]
port 410 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[16]
port 411 nsew signal input
rlabel metal3 s 119200 19048 120000 19168 6 la_oenb[17]
port 412 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 la_oenb[18]
port 413 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[19]
port 414 nsew signal input
rlabel metal3 s 119200 16328 120000 16448 6 la_oenb[1]
port 415 nsew signal input
rlabel metal3 s 119200 112208 120000 112328 6 la_oenb[20]
port 416 nsew signal input
rlabel metal3 s 119200 48968 120000 49088 6 la_oenb[21]
port 417 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[22]
port 418 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_oenb[23]
port 419 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[24]
port 420 nsew signal input
rlabel metal2 s 104990 119200 105046 120000 6 la_oenb[25]
port 421 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[26]
port 422 nsew signal input
rlabel metal3 s 119200 65288 120000 65408 6 la_oenb[27]
port 423 nsew signal input
rlabel metal2 s 119802 119200 119858 120000 6 la_oenb[28]
port 424 nsew signal input
rlabel metal2 s 106922 119200 106978 120000 6 la_oenb[29]
port 425 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 la_oenb[2]
port 426 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 la_oenb[30]
port 427 nsew signal input
rlabel metal2 s 35438 119200 35494 120000 6 la_oenb[31]
port 428 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_oenb[32]
port 429 nsew signal input
rlabel metal2 s 15474 119200 15530 120000 6 la_oenb[33]
port 430 nsew signal input
rlabel metal3 s 119200 37408 120000 37528 6 la_oenb[34]
port 431 nsew signal input
rlabel metal3 s 119200 69368 120000 69488 6 la_oenb[35]
port 432 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[36]
port 433 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[37]
port 434 nsew signal input
rlabel metal3 s 119200 97928 120000 98048 6 la_oenb[38]
port 435 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 la_oenb[39]
port 436 nsew signal input
rlabel metal2 s 109498 119200 109554 120000 6 la_oenb[3]
port 437 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 la_oenb[40]
port 438 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_oenb[41]
port 439 nsew signal input
rlabel metal2 s 7746 119200 7802 120000 6 la_oenb[42]
port 440 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 la_oenb[43]
port 441 nsew signal input
rlabel metal3 s 119200 5448 120000 5568 6 la_oenb[44]
port 442 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_oenb[45]
port 443 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_oenb[46]
port 444 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_oenb[47]
port 445 nsew signal input
rlabel metal3 s 119200 34688 120000 34808 6 la_oenb[48]
port 446 nsew signal input
rlabel metal3 s 119200 98608 120000 98728 6 la_oenb[49]
port 447 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 la_oenb[4]
port 448 nsew signal input
rlabel metal2 s 57334 119200 57390 120000 6 la_oenb[50]
port 449 nsew signal input
rlabel metal2 s 38658 119200 38714 120000 6 la_oenb[51]
port 450 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 la_oenb[52]
port 451 nsew signal input
rlabel metal3 s 119200 110848 120000 110968 6 la_oenb[53]
port 452 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 la_oenb[54]
port 453 nsew signal input
rlabel metal2 s 31574 119200 31630 120000 6 la_oenb[55]
port 454 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_oenb[56]
port 455 nsew signal input
rlabel metal3 s 119200 96568 120000 96688 6 la_oenb[57]
port 456 nsew signal input
rlabel metal2 s 84382 119200 84438 120000 6 la_oenb[58]
port 457 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 la_oenb[59]
port 458 nsew signal input
rlabel metal2 s 97262 119200 97318 120000 6 la_oenb[5]
port 459 nsew signal input
rlabel metal2 s 103702 119200 103758 120000 6 la_oenb[60]
port 460 nsew signal input
rlabel metal2 s 104346 119200 104402 120000 6 la_oenb[61]
port 461 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[62]
port 462 nsew signal input
rlabel metal2 s 65062 119200 65118 120000 6 la_oenb[63]
port 463 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_oenb[64]
port 464 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la_oenb[65]
port 465 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[66]
port 466 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 la_oenb[67]
port 467 nsew signal input
rlabel metal3 s 119200 22448 120000 22568 6 la_oenb[68]
port 468 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 la_oenb[69]
port 469 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 la_oenb[6]
port 470 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 la_oenb[70]
port 471 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_oenb[71]
port 472 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_oenb[72]
port 473 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la_oenb[73]
port 474 nsew signal input
rlabel metal2 s 61842 119200 61898 120000 6 la_oenb[74]
port 475 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[75]
port 476 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[76]
port 477 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 la_oenb[77]
port 478 nsew signal input
rlabel metal3 s 119200 82968 120000 83088 6 la_oenb[78]
port 479 nsew signal input
rlabel metal3 s 119200 108808 120000 108928 6 la_oenb[79]
port 480 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 la_oenb[7]
port 481 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 la_oenb[80]
port 482 nsew signal input
rlabel metal3 s 119200 12248 120000 12368 6 la_oenb[81]
port 483 nsew signal input
rlabel metal3 s 119200 102688 120000 102808 6 la_oenb[82]
port 484 nsew signal input
rlabel metal2 s 45742 119200 45798 120000 6 la_oenb[83]
port 485 nsew signal input
rlabel metal3 s 119200 85688 120000 85808 6 la_oenb[84]
port 486 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[85]
port 487 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_oenb[86]
port 488 nsew signal input
rlabel metal3 s 119200 26528 120000 26648 6 la_oenb[87]
port 489 nsew signal input
rlabel metal2 s 36082 119200 36138 120000 6 la_oenb[88]
port 490 nsew signal input
rlabel metal3 s 119200 2048 120000 2168 6 la_oenb[89]
port 491 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 la_oenb[8]
port 492 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 la_oenb[90]
port 493 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 la_oenb[91]
port 494 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[92]
port 495 nsew signal input
rlabel metal3 s 119200 102008 120000 102128 6 la_oenb[93]
port 496 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_oenb[94]
port 497 nsew signal input
rlabel metal3 s 119200 4088 120000 4208 6 la_oenb[95]
port 498 nsew signal input
rlabel metal2 s 662 119200 718 120000 6 la_oenb[96]
port 499 nsew signal input
rlabel metal2 s 74722 119200 74778 120000 6 la_oenb[97]
port 500 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 la_oenb[98]
port 501 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_oenb[99]
port 502 nsew signal input
rlabel metal2 s 8390 119200 8446 120000 6 la_oenb[9]
port 503 nsew signal input
rlabel metal4 s 5528 2128 5848 117552 6 vccd1
port 504 nsew power bidirectional
rlabel metal4 s 36248 2128 36568 117552 6 vccd1
port 504 nsew power bidirectional
rlabel metal4 s 66968 2128 67288 117552 6 vccd1
port 504 nsew power bidirectional
rlabel metal4 s 97688 2128 98008 117552 6 vccd1
port 504 nsew power bidirectional
rlabel metal5 s 1056 6666 118912 6986 6 vccd1
port 504 nsew power bidirectional
rlabel metal5 s 1056 37302 118912 37622 6 vccd1
port 504 nsew power bidirectional
rlabel metal5 s 1056 67938 118912 68258 6 vccd1
port 504 nsew power bidirectional
rlabel metal5 s 1056 98574 118912 98894 6 vccd1
port 504 nsew power bidirectional
rlabel metal4 s 6188 2128 6508 117552 6 vssd1
port 505 nsew ground bidirectional
rlabel metal4 s 36908 2128 37228 117552 6 vssd1
port 505 nsew ground bidirectional
rlabel metal4 s 67628 2128 67948 117552 6 vssd1
port 505 nsew ground bidirectional
rlabel metal4 s 98348 2128 98668 117552 6 vssd1
port 505 nsew ground bidirectional
rlabel metal5 s 1056 7326 118912 7646 6 vssd1
port 505 nsew ground bidirectional
rlabel metal5 s 1056 37962 118912 38282 6 vssd1
port 505 nsew ground bidirectional
rlabel metal5 s 1056 68598 118912 68918 6 vssd1
port 505 nsew ground bidirectional
rlabel metal5 s 1056 99234 118912 99554 6 vssd1
port 505 nsew ground bidirectional
rlabel metal3 s 119200 34008 120000 34128 6 wb_clk_i
port 506 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 wb_rst_i
port 507 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 wbs_ack_o
port 508 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 wbs_adr_i[0]
port 509 nsew signal input
rlabel metal2 s 25778 119200 25834 120000 6 wbs_adr_i[10]
port 510 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 wbs_adr_i[11]
port 511 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[12]
port 512 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 wbs_adr_i[13]
port 513 nsew signal input
rlabel metal3 s 119200 108128 120000 108248 6 wbs_adr_i[14]
port 514 nsew signal input
rlabel metal3 s 119200 99968 120000 100088 6 wbs_adr_i[15]
port 515 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 wbs_adr_i[16]
port 516 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 wbs_adr_i[17]
port 517 nsew signal input
rlabel metal3 s 119200 50328 120000 50448 6 wbs_adr_i[18]
port 518 nsew signal input
rlabel metal3 s 119200 2728 120000 2848 6 wbs_adr_i[19]
port 519 nsew signal input
rlabel metal2 s 54114 119200 54170 120000 6 wbs_adr_i[1]
port 520 nsew signal input
rlabel metal2 s 90178 119200 90234 120000 6 wbs_adr_i[20]
port 521 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_adr_i[21]
port 522 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 wbs_adr_i[22]
port 523 nsew signal input
rlabel metal3 s 119200 38088 120000 38208 6 wbs_adr_i[23]
port 524 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 wbs_adr_i[24]
port 525 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_adr_i[25]
port 526 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[26]
port 527 nsew signal input
rlabel metal2 s 18050 119200 18106 120000 6 wbs_adr_i[27]
port 528 nsew signal input
rlabel metal3 s 119200 83648 120000 83768 6 wbs_adr_i[28]
port 529 nsew signal input
rlabel metal2 s 107566 119200 107622 120000 6 wbs_adr_i[29]
port 530 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_adr_i[2]
port 531 nsew signal input
rlabel metal2 s 76654 119200 76710 120000 6 wbs_adr_i[30]
port 532 nsew signal input
rlabel metal3 s 119200 61888 120000 62008 6 wbs_adr_i[31]
port 533 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 wbs_adr_i[3]
port 534 nsew signal input
rlabel metal2 s 74078 119200 74134 120000 6 wbs_adr_i[4]
port 535 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 wbs_adr_i[5]
port 536 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_adr_i[6]
port 537 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[7]
port 538 nsew signal input
rlabel metal3 s 119200 4768 120000 4888 6 wbs_adr_i[8]
port 539 nsew signal input
rlabel metal3 s 119200 40808 120000 40928 6 wbs_adr_i[9]
port 540 nsew signal input
rlabel metal2 s 19338 119200 19394 120000 6 wbs_cyc_i
port 541 nsew signal input
rlabel metal3 s 119200 119688 120000 119808 6 wbs_dat_i[0]
port 542 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 wbs_dat_i[10]
port 543 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 wbs_dat_i[11]
port 544 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_dat_i[12]
port 545 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_dat_i[13]
port 546 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[14]
port 547 nsew signal input
rlabel metal3 s 119200 72088 120000 72208 6 wbs_dat_i[15]
port 548 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_i[16]
port 549 nsew signal input
rlabel metal2 s 68282 119200 68338 120000 6 wbs_dat_i[17]
port 550 nsew signal input
rlabel metal2 s 97906 119200 97962 120000 6 wbs_dat_i[18]
port 551 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 wbs_dat_i[19]
port 552 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[1]
port 553 nsew signal input
rlabel metal3 s 119200 81608 120000 81728 6 wbs_dat_i[20]
port 554 nsew signal input
rlabel metal2 s 103058 119200 103114 120000 6 wbs_dat_i[21]
port 555 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 wbs_dat_i[22]
port 556 nsew signal input
rlabel metal3 s 119200 104048 120000 104168 6 wbs_dat_i[23]
port 557 nsew signal input
rlabel metal3 s 119200 44888 120000 45008 6 wbs_dat_i[24]
port 558 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wbs_dat_i[25]
port 559 nsew signal input
rlabel metal2 s 89534 119200 89590 120000 6 wbs_dat_i[26]
port 560 nsew signal input
rlabel metal2 s 16762 119200 16818 120000 6 wbs_dat_i[27]
port 561 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[28]
port 562 nsew signal input
rlabel metal3 s 119200 79568 120000 79688 6 wbs_dat_i[29]
port 563 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_i[2]
port 564 nsew signal input
rlabel metal3 s 119200 39448 120000 39568 6 wbs_dat_i[30]
port 565 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 wbs_dat_i[31]
port 566 nsew signal input
rlabel metal3 s 119200 6128 120000 6248 6 wbs_dat_i[3]
port 567 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[4]
port 568 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_dat_i[5]
port 569 nsew signal input
rlabel metal3 s 119200 57128 120000 57248 6 wbs_dat_i[6]
port 570 nsew signal input
rlabel metal2 s 87602 119200 87658 120000 6 wbs_dat_i[7]
port 571 nsew signal input
rlabel metal3 s 119200 115608 120000 115728 6 wbs_dat_i[8]
port 572 nsew signal input
rlabel metal3 s 119200 6808 120000 6928 6 wbs_dat_i[9]
port 573 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[0]
port 574 nsew signal output
rlabel metal3 s 119200 73448 120000 73568 6 wbs_dat_o[10]
port 575 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_o[11]
port 576 nsew signal output
rlabel metal3 s 119200 116968 120000 117088 6 wbs_dat_o[12]
port 577 nsew signal output
rlabel metal2 s 83738 119200 83794 120000 6 wbs_dat_o[13]
port 578 nsew signal output
rlabel metal3 s 119200 14288 120000 14408 6 wbs_dat_o[14]
port 579 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 wbs_dat_o[15]
port 580 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 wbs_dat_o[16]
port 581 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 wbs_dat_o[17]
port 582 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 wbs_dat_o[18]
port 583 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 584 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_o[1]
port 585 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 wbs_dat_o[20]
port 586 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 wbs_dat_o[21]
port 587 nsew signal output
rlabel metal2 s 29642 119200 29698 120000 6 wbs_dat_o[22]
port 588 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 wbs_dat_o[23]
port 589 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[24]
port 590 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[25]
port 591 nsew signal output
rlabel metal2 s 59266 119200 59322 120000 6 wbs_dat_o[26]
port 592 nsew signal output
rlabel metal2 s 32218 119200 32274 120000 6 wbs_dat_o[27]
port 593 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 wbs_dat_o[28]
port 594 nsew signal output
rlabel metal2 s 80518 119200 80574 120000 6 wbs_dat_o[29]
port 595 nsew signal output
rlabel metal3 s 119200 33328 120000 33448 6 wbs_dat_o[2]
port 596 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 wbs_dat_o[30]
port 597 nsew signal output
rlabel metal3 s 119200 94528 120000 94648 6 wbs_dat_o[31]
port 598 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[3]
port 599 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_o[4]
port 600 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 wbs_dat_o[5]
port 601 nsew signal output
rlabel metal3 s 119200 89768 120000 89888 6 wbs_dat_o[6]
port 602 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 wbs_dat_o[7]
port 603 nsew signal output
rlabel metal2 s 77942 119200 77998 120000 6 wbs_dat_o[8]
port 604 nsew signal output
rlabel metal2 s 77298 119200 77354 120000 6 wbs_dat_o[9]
port 605 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 wbs_sel_i[0]
port 606 nsew signal input
rlabel metal2 s 14186 119200 14242 120000 6 wbs_sel_i[1]
port 607 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 wbs_sel_i[2]
port 608 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_sel_i[3]
port 609 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wbs_stb_i
port 610 nsew signal input
rlabel metal3 s 119200 57808 120000 57928 6 wbs_we_i
port 611 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6899276
string GDS_FILE /home/marwan/spm_ip/openlane/spm/runs/2023-03-22-11-30-24/results/signoff/spm.magic.gds
string GDS_START 361952
<< end >>

